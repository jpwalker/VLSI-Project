



ENTITY counter IS
	PORT(data_pass : IN BIT;
			msg_rdy : OUT BIT);
END counter;