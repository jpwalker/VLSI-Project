-- decoder_bdy.vhd
-- Jean P. Walker
-- File contains the body of the decoder package.

package body DecoderParts is
end package body;
