//
// Verilog description for cell multiplier, 
// Tue May  7 23:30:42 2019
//
// LeonardoSpectrum Level 3, 2011a.4 
//


module multiplier ( A_15__4, A_15__3, A_15__2, A_15__1, A_15__0, A_14__4, 
                    A_14__3, A_14__2, A_14__1, A_14__0, A_13__4, A_13__3, 
                    A_13__2, A_13__1, A_13__0, A_12__4, A_12__3, A_12__2, 
                    A_12__1, A_12__0, A_11__4, A_11__3, A_11__2, A_11__1, 
                    A_11__0, A_10__4, A_10__3, A_10__2, A_10__1, A_10__0, A_9__4, 
                    A_9__3, A_9__2, A_9__1, A_9__0, A_8__4, A_8__3, A_8__2, 
                    A_8__1, A_8__0, A_7__4, A_7__3, A_7__2, A_7__1, A_7__0, 
                    A_6__4, A_6__3, A_6__2, A_6__1, A_6__0, A_5__4, A_5__3, 
                    A_5__2, A_5__1, A_5__0, A_4__4, A_4__3, A_4__2, A_4__1, 
                    A_4__0, A_3__4, A_3__3, A_3__2, A_3__1, A_3__0, A_2__4, 
                    A_2__3, A_2__2, A_2__1, A_2__0, A_1__4, A_1__3, A_1__2, 
                    A_1__1, A_1__0, A_0__4, A_0__3, A_0__2, A_0__1, A_0__0, 
                    B_15__4, B_15__3, B_15__2, B_15__1, B_15__0, B_14__4, 
                    B_14__3, B_14__2, B_14__1, B_14__0, B_13__4, B_13__3, 
                    B_13__2, B_13__1, B_13__0, B_12__4, B_12__3, B_12__2, 
                    B_12__1, B_12__0, B_11__4, B_11__3, B_11__2, B_11__1, 
                    B_11__0, B_10__4, B_10__3, B_10__2, B_10__1, B_10__0, B_9__4, 
                    B_9__3, B_9__2, B_9__1, B_9__0, B_8__4, B_8__3, B_8__2, 
                    B_8__1, B_8__0, B_7__4, B_7__3, B_7__2, B_7__1, B_7__0, 
                    B_6__4, B_6__3, B_6__2, B_6__1, B_6__0, B_5__4, B_5__3, 
                    B_5__2, B_5__1, B_5__0, B_4__4, B_4__3, B_4__2, B_4__1, 
                    B_4__0, B_3__4, B_3__3, B_3__2, B_3__1, B_3__0, B_2__4, 
                    B_2__3, B_2__2, B_2__1, B_2__0, B_1__4, B_1__3, B_1__2, 
                    B_1__1, B_1__0, B_0__4, B_0__3, B_0__2, B_0__1, B_0__0, 
                    C_15__4, C_15__3, C_15__2, C_15__1, C_15__0, C_14__4, 
                    C_14__3, C_14__2, C_14__1, C_14__0, C_13__4, C_13__3, 
                    C_13__2, C_13__1, C_13__0, C_12__4, C_12__3, C_12__2, 
                    C_12__1, C_12__0, C_11__4, C_11__3, C_11__2, C_11__1, 
                    C_11__0, C_10__4, C_10__3, C_10__2, C_10__1, C_10__0, C_9__4, 
                    C_9__3, C_9__2, C_9__1, C_9__0, C_8__4, C_8__3, C_8__2, 
                    C_8__1, C_8__0, C_7__4, C_7__3, C_7__2, C_7__1, C_7__0, 
                    C_6__4, C_6__3, C_6__2, C_6__1, C_6__0, C_5__4, C_5__3, 
                    C_5__2, C_5__1, C_5__0, C_4__4, C_4__3, C_4__2, C_4__1, 
                    C_4__0, C_3__4, C_3__3, C_3__2, C_3__1, C_3__0, C_2__4, 
                    C_2__3, C_2__2, C_2__1, C_2__0, C_1__4, C_1__3, C_1__2, 
                    C_1__1, C_1__0, C_0__4, C_0__3, C_0__2, C_0__1, C_0__0 ) ;

    input A_15__4 ;
    input A_15__3 ;
    input A_15__2 ;
    input A_15__1 ;
    input A_15__0 ;
    input A_14__4 ;
    input A_14__3 ;
    input A_14__2 ;
    input A_14__1 ;
    input A_14__0 ;
    input A_13__4 ;
    input A_13__3 ;
    input A_13__2 ;
    input A_13__1 ;
    input A_13__0 ;
    input A_12__4 ;
    input A_12__3 ;
    input A_12__2 ;
    input A_12__1 ;
    input A_12__0 ;
    input A_11__4 ;
    input A_11__3 ;
    input A_11__2 ;
    input A_11__1 ;
    input A_11__0 ;
    input A_10__4 ;
    input A_10__3 ;
    input A_10__2 ;
    input A_10__1 ;
    input A_10__0 ;
    input A_9__4 ;
    input A_9__3 ;
    input A_9__2 ;
    input A_9__1 ;
    input A_9__0 ;
    input A_8__4 ;
    input A_8__3 ;
    input A_8__2 ;
    input A_8__1 ;
    input A_8__0 ;
    input A_7__4 ;
    input A_7__3 ;
    input A_7__2 ;
    input A_7__1 ;
    input A_7__0 ;
    input A_6__4 ;
    input A_6__3 ;
    input A_6__2 ;
    input A_6__1 ;
    input A_6__0 ;
    input A_5__4 ;
    input A_5__3 ;
    input A_5__2 ;
    input A_5__1 ;
    input A_5__0 ;
    input A_4__4 ;
    input A_4__3 ;
    input A_4__2 ;
    input A_4__1 ;
    input A_4__0 ;
    input A_3__4 ;
    input A_3__3 ;
    input A_3__2 ;
    input A_3__1 ;
    input A_3__0 ;
    input A_2__4 ;
    input A_2__3 ;
    input A_2__2 ;
    input A_2__1 ;
    input A_2__0 ;
    input A_1__4 ;
    input A_1__3 ;
    input A_1__2 ;
    input A_1__1 ;
    input A_1__0 ;
    input A_0__4 ;
    input A_0__3 ;
    input A_0__2 ;
    input A_0__1 ;
    input A_0__0 ;
    input B_15__4 ;
    input B_15__3 ;
    input B_15__2 ;
    input B_15__1 ;
    input B_15__0 ;
    input B_14__4 ;
    input B_14__3 ;
    input B_14__2 ;
    input B_14__1 ;
    input B_14__0 ;
    input B_13__4 ;
    input B_13__3 ;
    input B_13__2 ;
    input B_13__1 ;
    input B_13__0 ;
    input B_12__4 ;
    input B_12__3 ;
    input B_12__2 ;
    input B_12__1 ;
    input B_12__0 ;
    input B_11__4 ;
    input B_11__3 ;
    input B_11__2 ;
    input B_11__1 ;
    input B_11__0 ;
    input B_10__4 ;
    input B_10__3 ;
    input B_10__2 ;
    input B_10__1 ;
    input B_10__0 ;
    input B_9__4 ;
    input B_9__3 ;
    input B_9__2 ;
    input B_9__1 ;
    input B_9__0 ;
    input B_8__4 ;
    input B_8__3 ;
    input B_8__2 ;
    input B_8__1 ;
    input B_8__0 ;
    input B_7__4 ;
    input B_7__3 ;
    input B_7__2 ;
    input B_7__1 ;
    input B_7__0 ;
    input B_6__4 ;
    input B_6__3 ;
    input B_6__2 ;
    input B_6__1 ;
    input B_6__0 ;
    input B_5__4 ;
    input B_5__3 ;
    input B_5__2 ;
    input B_5__1 ;
    input B_5__0 ;
    input B_4__4 ;
    input B_4__3 ;
    input B_4__2 ;
    input B_4__1 ;
    input B_4__0 ;
    input B_3__4 ;
    input B_3__3 ;
    input B_3__2 ;
    input B_3__1 ;
    input B_3__0 ;
    input B_2__4 ;
    input B_2__3 ;
    input B_2__2 ;
    input B_2__1 ;
    input B_2__0 ;
    input B_1__4 ;
    input B_1__3 ;
    input B_1__2 ;
    input B_1__1 ;
    input B_1__0 ;
    input B_0__4 ;
    input B_0__3 ;
    input B_0__2 ;
    input B_0__1 ;
    input B_0__0 ;
    output C_15__4 ;
    output C_15__3 ;
    output C_15__2 ;
    output C_15__1 ;
    output C_15__0 ;
    output C_14__4 ;
    output C_14__3 ;
    output C_14__2 ;
    output C_14__1 ;
    output C_14__0 ;
    output C_13__4 ;
    output C_13__3 ;
    output C_13__2 ;
    output C_13__1 ;
    output C_13__0 ;
    output C_12__4 ;
    output C_12__3 ;
    output C_12__2 ;
    output C_12__1 ;
    output C_12__0 ;
    output C_11__4 ;
    output C_11__3 ;
    output C_11__2 ;
    output C_11__1 ;
    output C_11__0 ;
    output C_10__4 ;
    output C_10__3 ;
    output C_10__2 ;
    output C_10__1 ;
    output C_10__0 ;
    output C_9__4 ;
    output C_9__3 ;
    output C_9__2 ;
    output C_9__1 ;
    output C_9__0 ;
    output C_8__4 ;
    output C_8__3 ;
    output C_8__2 ;
    output C_8__1 ;
    output C_8__0 ;
    output C_7__4 ;
    output C_7__3 ;
    output C_7__2 ;
    output C_7__1 ;
    output C_7__0 ;
    output C_6__4 ;
    output C_6__3 ;
    output C_6__2 ;
    output C_6__1 ;
    output C_6__0 ;
    output C_5__4 ;
    output C_5__3 ;
    output C_5__2 ;
    output C_5__1 ;
    output C_5__0 ;
    output C_4__4 ;
    output C_4__3 ;
    output C_4__2 ;
    output C_4__1 ;
    output C_4__0 ;
    output C_3__4 ;
    output C_3__3 ;
    output C_3__2 ;
    output C_3__1 ;
    output C_3__0 ;
    output C_2__4 ;
    output C_2__3 ;
    output C_2__2 ;
    output C_2__1 ;
    output C_2__0 ;
    output C_1__4 ;
    output C_1__3 ;
    output C_1__2 ;
    output C_1__1 ;
    output C_1__0 ;
    output C_0__4 ;
    output C_0__3 ;
    output C_0__2 ;
    output C_0__1 ;
    output C_0__0 ;

    wire chipmulties_15_cm_nx2, chipmulties_15_cm_nx10, chipmulties_15_cm_nx12, 
         chipmulties_15_cm_nx14, chipmulties_15_cm_nx18, chipmulties_15_cm_nx22, 
         chipmulties_15_cm_nx28, chipmulties_15_cm_nx46, chipmulties_15_cm_nx52, 
         chipmulties_15_cm_nx54, chipmulties_15_cm_nx62, chipmulties_15_cm_nx68, 
         chipmulties_15_cm_nx78, chipmulties_15_cm_nx118, 
         chipmulties_15_cm_nx130, chipmulties_15_cm_nx154, 
         chipmulties_15_cm_nx164, chipmulties_15_cm_nx178, 
         chipmulties_15_cm_nx192, chipmulties_15_cm_nx228, 
         chipmulties_15_cm_nx501, chipmulties_15_cm_nx503, 
         chipmulties_15_cm_nx506, chipmulties_15_cm_nx508, 
         chipmulties_15_cm_nx511, chipmulties_15_cm_nx513, 
         chipmulties_15_cm_nx518, chipmulties_15_cm_nx523, 
         chipmulties_15_cm_nx528, chipmulties_15_cm_nx533, 
         chipmulties_15_cm_nx535, chipmulties_15_cm_nx537, 
         chipmulties_15_cm_nx539, chipmulties_15_cm_nx541, 
         chipmulties_15_cm_nx543, chipmulties_15_cm_nx545, 
         chipmulties_15_cm_nx547, chipmulties_15_cm_nx550, 
         chipmulties_15_cm_nx553, chipmulties_15_cm_nx555, 
         chipmulties_15_cm_nx557, chipmulties_15_cm_nx560, 
         chipmulties_15_cm_nx562, chipmulties_15_cm_nx566, 
         chipmulties_15_cm_nx569, chipmulties_15_cm_nx571, 
         chipmulties_15_cm_nx573, chipmulties_15_cm_nx575, 
         chipmulties_15_cm_nx580, chipmulties_15_cm_nx583, 
         chipmulties_15_cm_nx587, chipmulties_15_cm_nx589, 
         chipmulties_15_cm_nx591, chipmulties_14_cm_nx2, chipmulties_14_cm_nx10, 
         chipmulties_14_cm_nx12, chipmulties_14_cm_nx14, chipmulties_14_cm_nx18, 
         chipmulties_14_cm_nx22, chipmulties_14_cm_nx28, chipmulties_14_cm_nx46, 
         chipmulties_14_cm_nx52, chipmulties_14_cm_nx54, chipmulties_14_cm_nx62, 
         chipmulties_14_cm_nx68, chipmulties_14_cm_nx78, chipmulties_14_cm_nx118, 
         chipmulties_14_cm_nx130, chipmulties_14_cm_nx154, 
         chipmulties_14_cm_nx164, chipmulties_14_cm_nx178, 
         chipmulties_14_cm_nx192, chipmulties_14_cm_nx228, 
         chipmulties_14_cm_nx501, chipmulties_14_cm_nx503, 
         chipmulties_14_cm_nx506, chipmulties_14_cm_nx508, 
         chipmulties_14_cm_nx511, chipmulties_14_cm_nx513, 
         chipmulties_14_cm_nx518, chipmulties_14_cm_nx523, 
         chipmulties_14_cm_nx528, chipmulties_14_cm_nx533, 
         chipmulties_14_cm_nx535, chipmulties_14_cm_nx537, 
         chipmulties_14_cm_nx539, chipmulties_14_cm_nx541, 
         chipmulties_14_cm_nx543, chipmulties_14_cm_nx545, 
         chipmulties_14_cm_nx547, chipmulties_14_cm_nx550, 
         chipmulties_14_cm_nx553, chipmulties_14_cm_nx555, 
         chipmulties_14_cm_nx557, chipmulties_14_cm_nx560, 
         chipmulties_14_cm_nx562, chipmulties_14_cm_nx566, 
         chipmulties_14_cm_nx569, chipmulties_14_cm_nx571, 
         chipmulties_14_cm_nx573, chipmulties_14_cm_nx575, 
         chipmulties_14_cm_nx580, chipmulties_14_cm_nx583, 
         chipmulties_14_cm_nx587, chipmulties_14_cm_nx589, 
         chipmulties_14_cm_nx591, chipmulties_13_cm_nx2, chipmulties_13_cm_nx10, 
         chipmulties_13_cm_nx12, chipmulties_13_cm_nx14, chipmulties_13_cm_nx18, 
         chipmulties_13_cm_nx22, chipmulties_13_cm_nx28, chipmulties_13_cm_nx46, 
         chipmulties_13_cm_nx52, chipmulties_13_cm_nx54, chipmulties_13_cm_nx62, 
         chipmulties_13_cm_nx68, chipmulties_13_cm_nx78, chipmulties_13_cm_nx118, 
         chipmulties_13_cm_nx130, chipmulties_13_cm_nx154, 
         chipmulties_13_cm_nx164, chipmulties_13_cm_nx178, 
         chipmulties_13_cm_nx192, chipmulties_13_cm_nx228, 
         chipmulties_13_cm_nx501, chipmulties_13_cm_nx503, 
         chipmulties_13_cm_nx506, chipmulties_13_cm_nx508, 
         chipmulties_13_cm_nx511, chipmulties_13_cm_nx513, 
         chipmulties_13_cm_nx518, chipmulties_13_cm_nx523, 
         chipmulties_13_cm_nx528, chipmulties_13_cm_nx533, 
         chipmulties_13_cm_nx535, chipmulties_13_cm_nx537, 
         chipmulties_13_cm_nx539, chipmulties_13_cm_nx541, 
         chipmulties_13_cm_nx543, chipmulties_13_cm_nx545, 
         chipmulties_13_cm_nx547, chipmulties_13_cm_nx550, 
         chipmulties_13_cm_nx553, chipmulties_13_cm_nx555, 
         chipmulties_13_cm_nx557, chipmulties_13_cm_nx560, 
         chipmulties_13_cm_nx562, chipmulties_13_cm_nx566, 
         chipmulties_13_cm_nx569, chipmulties_13_cm_nx571, 
         chipmulties_13_cm_nx573, chipmulties_13_cm_nx575, 
         chipmulties_13_cm_nx580, chipmulties_13_cm_nx583, 
         chipmulties_13_cm_nx587, chipmulties_13_cm_nx589, 
         chipmulties_13_cm_nx591, chipmulties_12_cm_nx2, chipmulties_12_cm_nx10, 
         chipmulties_12_cm_nx12, chipmulties_12_cm_nx14, chipmulties_12_cm_nx18, 
         chipmulties_12_cm_nx22, chipmulties_12_cm_nx28, chipmulties_12_cm_nx46, 
         chipmulties_12_cm_nx52, chipmulties_12_cm_nx54, chipmulties_12_cm_nx62, 
         chipmulties_12_cm_nx68, chipmulties_12_cm_nx78, chipmulties_12_cm_nx118, 
         chipmulties_12_cm_nx130, chipmulties_12_cm_nx154, 
         chipmulties_12_cm_nx164, chipmulties_12_cm_nx178, 
         chipmulties_12_cm_nx192, chipmulties_12_cm_nx228, 
         chipmulties_12_cm_nx501, chipmulties_12_cm_nx503, 
         chipmulties_12_cm_nx506, chipmulties_12_cm_nx508, 
         chipmulties_12_cm_nx511, chipmulties_12_cm_nx513, 
         chipmulties_12_cm_nx518, chipmulties_12_cm_nx523, 
         chipmulties_12_cm_nx528, chipmulties_12_cm_nx533, 
         chipmulties_12_cm_nx535, chipmulties_12_cm_nx537, 
         chipmulties_12_cm_nx539, chipmulties_12_cm_nx541, 
         chipmulties_12_cm_nx543, chipmulties_12_cm_nx545, 
         chipmulties_12_cm_nx547, chipmulties_12_cm_nx550, 
         chipmulties_12_cm_nx553, chipmulties_12_cm_nx555, 
         chipmulties_12_cm_nx557, chipmulties_12_cm_nx560, 
         chipmulties_12_cm_nx562, chipmulties_12_cm_nx566, 
         chipmulties_12_cm_nx569, chipmulties_12_cm_nx571, 
         chipmulties_12_cm_nx573, chipmulties_12_cm_nx575, 
         chipmulties_12_cm_nx580, chipmulties_12_cm_nx583, 
         chipmulties_12_cm_nx587, chipmulties_12_cm_nx589, 
         chipmulties_12_cm_nx591, chipmulties_11_cm_nx2, chipmulties_11_cm_nx10, 
         chipmulties_11_cm_nx12, chipmulties_11_cm_nx14, chipmulties_11_cm_nx18, 
         chipmulties_11_cm_nx22, chipmulties_11_cm_nx28, chipmulties_11_cm_nx46, 
         chipmulties_11_cm_nx52, chipmulties_11_cm_nx54, chipmulties_11_cm_nx62, 
         chipmulties_11_cm_nx68, chipmulties_11_cm_nx78, chipmulties_11_cm_nx118, 
         chipmulties_11_cm_nx130, chipmulties_11_cm_nx154, 
         chipmulties_11_cm_nx164, chipmulties_11_cm_nx178, 
         chipmulties_11_cm_nx192, chipmulties_11_cm_nx228, 
         chipmulties_11_cm_nx501, chipmulties_11_cm_nx503, 
         chipmulties_11_cm_nx506, chipmulties_11_cm_nx508, 
         chipmulties_11_cm_nx511, chipmulties_11_cm_nx513, 
         chipmulties_11_cm_nx518, chipmulties_11_cm_nx523, 
         chipmulties_11_cm_nx528, chipmulties_11_cm_nx533, 
         chipmulties_11_cm_nx535, chipmulties_11_cm_nx537, 
         chipmulties_11_cm_nx539, chipmulties_11_cm_nx541, 
         chipmulties_11_cm_nx543, chipmulties_11_cm_nx545, 
         chipmulties_11_cm_nx547, chipmulties_11_cm_nx550, 
         chipmulties_11_cm_nx553, chipmulties_11_cm_nx555, 
         chipmulties_11_cm_nx557, chipmulties_11_cm_nx560, 
         chipmulties_11_cm_nx562, chipmulties_11_cm_nx566, 
         chipmulties_11_cm_nx569, chipmulties_11_cm_nx571, 
         chipmulties_11_cm_nx573, chipmulties_11_cm_nx575, 
         chipmulties_11_cm_nx580, chipmulties_11_cm_nx583, 
         chipmulties_11_cm_nx587, chipmulties_11_cm_nx589, 
         chipmulties_11_cm_nx591, chipmulties_10_cm_nx2, chipmulties_10_cm_nx10, 
         chipmulties_10_cm_nx12, chipmulties_10_cm_nx14, chipmulties_10_cm_nx18, 
         chipmulties_10_cm_nx22, chipmulties_10_cm_nx28, chipmulties_10_cm_nx46, 
         chipmulties_10_cm_nx52, chipmulties_10_cm_nx54, chipmulties_10_cm_nx62, 
         chipmulties_10_cm_nx68, chipmulties_10_cm_nx78, chipmulties_10_cm_nx118, 
         chipmulties_10_cm_nx130, chipmulties_10_cm_nx154, 
         chipmulties_10_cm_nx164, chipmulties_10_cm_nx178, 
         chipmulties_10_cm_nx192, chipmulties_10_cm_nx228, 
         chipmulties_10_cm_nx501, chipmulties_10_cm_nx503, 
         chipmulties_10_cm_nx506, chipmulties_10_cm_nx508, 
         chipmulties_10_cm_nx511, chipmulties_10_cm_nx513, 
         chipmulties_10_cm_nx518, chipmulties_10_cm_nx523, 
         chipmulties_10_cm_nx528, chipmulties_10_cm_nx533, 
         chipmulties_10_cm_nx535, chipmulties_10_cm_nx537, 
         chipmulties_10_cm_nx539, chipmulties_10_cm_nx541, 
         chipmulties_10_cm_nx543, chipmulties_10_cm_nx545, 
         chipmulties_10_cm_nx547, chipmulties_10_cm_nx550, 
         chipmulties_10_cm_nx553, chipmulties_10_cm_nx555, 
         chipmulties_10_cm_nx557, chipmulties_10_cm_nx560, 
         chipmulties_10_cm_nx562, chipmulties_10_cm_nx566, 
         chipmulties_10_cm_nx569, chipmulties_10_cm_nx571, 
         chipmulties_10_cm_nx573, chipmulties_10_cm_nx575, 
         chipmulties_10_cm_nx580, chipmulties_10_cm_nx583, 
         chipmulties_10_cm_nx587, chipmulties_10_cm_nx589, 
         chipmulties_10_cm_nx591, chipmulties_9_cm_nx2, chipmulties_9_cm_nx10, 
         chipmulties_9_cm_nx12, chipmulties_9_cm_nx14, chipmulties_9_cm_nx18, 
         chipmulties_9_cm_nx22, chipmulties_9_cm_nx28, chipmulties_9_cm_nx46, 
         chipmulties_9_cm_nx52, chipmulties_9_cm_nx54, chipmulties_9_cm_nx62, 
         chipmulties_9_cm_nx68, chipmulties_9_cm_nx78, chipmulties_9_cm_nx118, 
         chipmulties_9_cm_nx130, chipmulties_9_cm_nx154, chipmulties_9_cm_nx164, 
         chipmulties_9_cm_nx178, chipmulties_9_cm_nx192, chipmulties_9_cm_nx228, 
         chipmulties_9_cm_nx501, chipmulties_9_cm_nx503, chipmulties_9_cm_nx506, 
         chipmulties_9_cm_nx508, chipmulties_9_cm_nx511, chipmulties_9_cm_nx513, 
         chipmulties_9_cm_nx518, chipmulties_9_cm_nx523, chipmulties_9_cm_nx528, 
         chipmulties_9_cm_nx533, chipmulties_9_cm_nx535, chipmulties_9_cm_nx537, 
         chipmulties_9_cm_nx539, chipmulties_9_cm_nx541, chipmulties_9_cm_nx543, 
         chipmulties_9_cm_nx545, chipmulties_9_cm_nx547, chipmulties_9_cm_nx550, 
         chipmulties_9_cm_nx553, chipmulties_9_cm_nx555, chipmulties_9_cm_nx557, 
         chipmulties_9_cm_nx560, chipmulties_9_cm_nx562, chipmulties_9_cm_nx566, 
         chipmulties_9_cm_nx569, chipmulties_9_cm_nx571, chipmulties_9_cm_nx573, 
         chipmulties_9_cm_nx575, chipmulties_9_cm_nx580, chipmulties_9_cm_nx583, 
         chipmulties_9_cm_nx587, chipmulties_9_cm_nx589, chipmulties_9_cm_nx591, 
         chipmulties_8_cm_nx2, chipmulties_8_cm_nx10, chipmulties_8_cm_nx12, 
         chipmulties_8_cm_nx14, chipmulties_8_cm_nx18, chipmulties_8_cm_nx22, 
         chipmulties_8_cm_nx28, chipmulties_8_cm_nx46, chipmulties_8_cm_nx52, 
         chipmulties_8_cm_nx54, chipmulties_8_cm_nx62, chipmulties_8_cm_nx68, 
         chipmulties_8_cm_nx78, chipmulties_8_cm_nx118, chipmulties_8_cm_nx130, 
         chipmulties_8_cm_nx154, chipmulties_8_cm_nx164, chipmulties_8_cm_nx178, 
         chipmulties_8_cm_nx192, chipmulties_8_cm_nx228, chipmulties_8_cm_nx501, 
         chipmulties_8_cm_nx503, chipmulties_8_cm_nx506, chipmulties_8_cm_nx508, 
         chipmulties_8_cm_nx511, chipmulties_8_cm_nx513, chipmulties_8_cm_nx518, 
         chipmulties_8_cm_nx523, chipmulties_8_cm_nx528, chipmulties_8_cm_nx533, 
         chipmulties_8_cm_nx535, chipmulties_8_cm_nx537, chipmulties_8_cm_nx539, 
         chipmulties_8_cm_nx541, chipmulties_8_cm_nx543, chipmulties_8_cm_nx545, 
         chipmulties_8_cm_nx547, chipmulties_8_cm_nx550, chipmulties_8_cm_nx553, 
         chipmulties_8_cm_nx555, chipmulties_8_cm_nx557, chipmulties_8_cm_nx560, 
         chipmulties_8_cm_nx562, chipmulties_8_cm_nx566, chipmulties_8_cm_nx569, 
         chipmulties_8_cm_nx571, chipmulties_8_cm_nx573, chipmulties_8_cm_nx575, 
         chipmulties_8_cm_nx580, chipmulties_8_cm_nx583, chipmulties_8_cm_nx587, 
         chipmulties_8_cm_nx589, chipmulties_8_cm_nx591, chipmulties_7_cm_nx2, 
         chipmulties_7_cm_nx10, chipmulties_7_cm_nx12, chipmulties_7_cm_nx14, 
         chipmulties_7_cm_nx18, chipmulties_7_cm_nx22, chipmulties_7_cm_nx28, 
         chipmulties_7_cm_nx46, chipmulties_7_cm_nx52, chipmulties_7_cm_nx54, 
         chipmulties_7_cm_nx62, chipmulties_7_cm_nx68, chipmulties_7_cm_nx78, 
         chipmulties_7_cm_nx118, chipmulties_7_cm_nx130, chipmulties_7_cm_nx154, 
         chipmulties_7_cm_nx164, chipmulties_7_cm_nx178, chipmulties_7_cm_nx192, 
         chipmulties_7_cm_nx228, chipmulties_7_cm_nx501, chipmulties_7_cm_nx503, 
         chipmulties_7_cm_nx506, chipmulties_7_cm_nx508, chipmulties_7_cm_nx511, 
         chipmulties_7_cm_nx513, chipmulties_7_cm_nx518, chipmulties_7_cm_nx523, 
         chipmulties_7_cm_nx528, chipmulties_7_cm_nx533, chipmulties_7_cm_nx535, 
         chipmulties_7_cm_nx537, chipmulties_7_cm_nx539, chipmulties_7_cm_nx541, 
         chipmulties_7_cm_nx543, chipmulties_7_cm_nx545, chipmulties_7_cm_nx547, 
         chipmulties_7_cm_nx550, chipmulties_7_cm_nx553, chipmulties_7_cm_nx555, 
         chipmulties_7_cm_nx557, chipmulties_7_cm_nx560, chipmulties_7_cm_nx562, 
         chipmulties_7_cm_nx566, chipmulties_7_cm_nx569, chipmulties_7_cm_nx571, 
         chipmulties_7_cm_nx573, chipmulties_7_cm_nx575, chipmulties_7_cm_nx580, 
         chipmulties_7_cm_nx583, chipmulties_7_cm_nx587, chipmulties_7_cm_nx589, 
         chipmulties_7_cm_nx591, chipmulties_6_cm_nx2, chipmulties_6_cm_nx10, 
         chipmulties_6_cm_nx12, chipmulties_6_cm_nx14, chipmulties_6_cm_nx18, 
         chipmulties_6_cm_nx22, chipmulties_6_cm_nx28, chipmulties_6_cm_nx46, 
         chipmulties_6_cm_nx52, chipmulties_6_cm_nx54, chipmulties_6_cm_nx62, 
         chipmulties_6_cm_nx68, chipmulties_6_cm_nx78, chipmulties_6_cm_nx118, 
         chipmulties_6_cm_nx130, chipmulties_6_cm_nx154, chipmulties_6_cm_nx164, 
         chipmulties_6_cm_nx178, chipmulties_6_cm_nx192, chipmulties_6_cm_nx228, 
         chipmulties_6_cm_nx501, chipmulties_6_cm_nx503, chipmulties_6_cm_nx506, 
         chipmulties_6_cm_nx508, chipmulties_6_cm_nx511, chipmulties_6_cm_nx513, 
         chipmulties_6_cm_nx518, chipmulties_6_cm_nx523, chipmulties_6_cm_nx528, 
         chipmulties_6_cm_nx533, chipmulties_6_cm_nx535, chipmulties_6_cm_nx537, 
         chipmulties_6_cm_nx539, chipmulties_6_cm_nx541, chipmulties_6_cm_nx543, 
         chipmulties_6_cm_nx545, chipmulties_6_cm_nx547, chipmulties_6_cm_nx550, 
         chipmulties_6_cm_nx553, chipmulties_6_cm_nx555, chipmulties_6_cm_nx557, 
         chipmulties_6_cm_nx560, chipmulties_6_cm_nx562, chipmulties_6_cm_nx566, 
         chipmulties_6_cm_nx569, chipmulties_6_cm_nx571, chipmulties_6_cm_nx573, 
         chipmulties_6_cm_nx575, chipmulties_6_cm_nx580, chipmulties_6_cm_nx583, 
         chipmulties_6_cm_nx587, chipmulties_6_cm_nx589, chipmulties_6_cm_nx591, 
         chipmulties_5_cm_nx2, chipmulties_5_cm_nx10, chipmulties_5_cm_nx12, 
         chipmulties_5_cm_nx14, chipmulties_5_cm_nx18, chipmulties_5_cm_nx22, 
         chipmulties_5_cm_nx28, chipmulties_5_cm_nx46, chipmulties_5_cm_nx52, 
         chipmulties_5_cm_nx54, chipmulties_5_cm_nx62, chipmulties_5_cm_nx68, 
         chipmulties_5_cm_nx78, chipmulties_5_cm_nx118, chipmulties_5_cm_nx130, 
         chipmulties_5_cm_nx154, chipmulties_5_cm_nx164, chipmulties_5_cm_nx178, 
         chipmulties_5_cm_nx192, chipmulties_5_cm_nx228, chipmulties_5_cm_nx501, 
         chipmulties_5_cm_nx503, chipmulties_5_cm_nx506, chipmulties_5_cm_nx508, 
         chipmulties_5_cm_nx511, chipmulties_5_cm_nx513, chipmulties_5_cm_nx518, 
         chipmulties_5_cm_nx523, chipmulties_5_cm_nx528, chipmulties_5_cm_nx533, 
         chipmulties_5_cm_nx535, chipmulties_5_cm_nx537, chipmulties_5_cm_nx539, 
         chipmulties_5_cm_nx541, chipmulties_5_cm_nx543, chipmulties_5_cm_nx545, 
         chipmulties_5_cm_nx547, chipmulties_5_cm_nx550, chipmulties_5_cm_nx553, 
         chipmulties_5_cm_nx555, chipmulties_5_cm_nx557, chipmulties_5_cm_nx560, 
         chipmulties_5_cm_nx562, chipmulties_5_cm_nx566, chipmulties_5_cm_nx569, 
         chipmulties_5_cm_nx571, chipmulties_5_cm_nx573, chipmulties_5_cm_nx575, 
         chipmulties_5_cm_nx580, chipmulties_5_cm_nx583, chipmulties_5_cm_nx587, 
         chipmulties_5_cm_nx589, chipmulties_5_cm_nx591, chipmulties_4_cm_nx2, 
         chipmulties_4_cm_nx10, chipmulties_4_cm_nx12, chipmulties_4_cm_nx14, 
         chipmulties_4_cm_nx18, chipmulties_4_cm_nx22, chipmulties_4_cm_nx28, 
         chipmulties_4_cm_nx46, chipmulties_4_cm_nx52, chipmulties_4_cm_nx54, 
         chipmulties_4_cm_nx62, chipmulties_4_cm_nx68, chipmulties_4_cm_nx78, 
         chipmulties_4_cm_nx118, chipmulties_4_cm_nx130, chipmulties_4_cm_nx154, 
         chipmulties_4_cm_nx164, chipmulties_4_cm_nx178, chipmulties_4_cm_nx192, 
         chipmulties_4_cm_nx228, chipmulties_4_cm_nx501, chipmulties_4_cm_nx503, 
         chipmulties_4_cm_nx506, chipmulties_4_cm_nx508, chipmulties_4_cm_nx511, 
         chipmulties_4_cm_nx513, chipmulties_4_cm_nx518, chipmulties_4_cm_nx523, 
         chipmulties_4_cm_nx528, chipmulties_4_cm_nx533, chipmulties_4_cm_nx535, 
         chipmulties_4_cm_nx537, chipmulties_4_cm_nx539, chipmulties_4_cm_nx541, 
         chipmulties_4_cm_nx543, chipmulties_4_cm_nx545, chipmulties_4_cm_nx547, 
         chipmulties_4_cm_nx550, chipmulties_4_cm_nx553, chipmulties_4_cm_nx555, 
         chipmulties_4_cm_nx557, chipmulties_4_cm_nx560, chipmulties_4_cm_nx562, 
         chipmulties_4_cm_nx566, chipmulties_4_cm_nx569, chipmulties_4_cm_nx571, 
         chipmulties_4_cm_nx573, chipmulties_4_cm_nx575, chipmulties_4_cm_nx580, 
         chipmulties_4_cm_nx583, chipmulties_4_cm_nx587, chipmulties_4_cm_nx589, 
         chipmulties_4_cm_nx591, chipmulties_3_cm_nx2, chipmulties_3_cm_nx10, 
         chipmulties_3_cm_nx12, chipmulties_3_cm_nx14, chipmulties_3_cm_nx18, 
         chipmulties_3_cm_nx22, chipmulties_3_cm_nx28, chipmulties_3_cm_nx46, 
         chipmulties_3_cm_nx52, chipmulties_3_cm_nx54, chipmulties_3_cm_nx62, 
         chipmulties_3_cm_nx68, chipmulties_3_cm_nx78, chipmulties_3_cm_nx118, 
         chipmulties_3_cm_nx130, chipmulties_3_cm_nx154, chipmulties_3_cm_nx164, 
         chipmulties_3_cm_nx178, chipmulties_3_cm_nx192, chipmulties_3_cm_nx228, 
         chipmulties_3_cm_nx501, chipmulties_3_cm_nx503, chipmulties_3_cm_nx506, 
         chipmulties_3_cm_nx508, chipmulties_3_cm_nx511, chipmulties_3_cm_nx513, 
         chipmulties_3_cm_nx518, chipmulties_3_cm_nx523, chipmulties_3_cm_nx528, 
         chipmulties_3_cm_nx533, chipmulties_3_cm_nx535, chipmulties_3_cm_nx537, 
         chipmulties_3_cm_nx539, chipmulties_3_cm_nx541, chipmulties_3_cm_nx543, 
         chipmulties_3_cm_nx545, chipmulties_3_cm_nx547, chipmulties_3_cm_nx550, 
         chipmulties_3_cm_nx553, chipmulties_3_cm_nx555, chipmulties_3_cm_nx557, 
         chipmulties_3_cm_nx560, chipmulties_3_cm_nx562, chipmulties_3_cm_nx566, 
         chipmulties_3_cm_nx569, chipmulties_3_cm_nx571, chipmulties_3_cm_nx573, 
         chipmulties_3_cm_nx575, chipmulties_3_cm_nx580, chipmulties_3_cm_nx583, 
         chipmulties_3_cm_nx587, chipmulties_3_cm_nx589, chipmulties_3_cm_nx591, 
         chipmulties_2_cm_nx2, chipmulties_2_cm_nx10, chipmulties_2_cm_nx12, 
         chipmulties_2_cm_nx14, chipmulties_2_cm_nx18, chipmulties_2_cm_nx22, 
         chipmulties_2_cm_nx28, chipmulties_2_cm_nx46, chipmulties_2_cm_nx52, 
         chipmulties_2_cm_nx54, chipmulties_2_cm_nx62, chipmulties_2_cm_nx68, 
         chipmulties_2_cm_nx78, chipmulties_2_cm_nx118, chipmulties_2_cm_nx130, 
         chipmulties_2_cm_nx154, chipmulties_2_cm_nx164, chipmulties_2_cm_nx178, 
         chipmulties_2_cm_nx192, chipmulties_2_cm_nx228, chipmulties_2_cm_nx501, 
         chipmulties_2_cm_nx503, chipmulties_2_cm_nx506, chipmulties_2_cm_nx508, 
         chipmulties_2_cm_nx511, chipmulties_2_cm_nx513, chipmulties_2_cm_nx518, 
         chipmulties_2_cm_nx523, chipmulties_2_cm_nx528, chipmulties_2_cm_nx533, 
         chipmulties_2_cm_nx535, chipmulties_2_cm_nx537, chipmulties_2_cm_nx539, 
         chipmulties_2_cm_nx541, chipmulties_2_cm_nx543, chipmulties_2_cm_nx545, 
         chipmulties_2_cm_nx547, chipmulties_2_cm_nx550, chipmulties_2_cm_nx553, 
         chipmulties_2_cm_nx555, chipmulties_2_cm_nx557, chipmulties_2_cm_nx560, 
         chipmulties_2_cm_nx562, chipmulties_2_cm_nx566, chipmulties_2_cm_nx569, 
         chipmulties_2_cm_nx571, chipmulties_2_cm_nx573, chipmulties_2_cm_nx575, 
         chipmulties_2_cm_nx580, chipmulties_2_cm_nx583, chipmulties_2_cm_nx587, 
         chipmulties_2_cm_nx589, chipmulties_2_cm_nx591, chipmulties_1_cm_nx2, 
         chipmulties_1_cm_nx10, chipmulties_1_cm_nx12, chipmulties_1_cm_nx14, 
         chipmulties_1_cm_nx18, chipmulties_1_cm_nx22, chipmulties_1_cm_nx28, 
         chipmulties_1_cm_nx46, chipmulties_1_cm_nx52, chipmulties_1_cm_nx54, 
         chipmulties_1_cm_nx62, chipmulties_1_cm_nx68, chipmulties_1_cm_nx78, 
         chipmulties_1_cm_nx118, chipmulties_1_cm_nx130, chipmulties_1_cm_nx154, 
         chipmulties_1_cm_nx164, chipmulties_1_cm_nx178, chipmulties_1_cm_nx192, 
         chipmulties_1_cm_nx228, chipmulties_1_cm_nx501, chipmulties_1_cm_nx503, 
         chipmulties_1_cm_nx506, chipmulties_1_cm_nx508, chipmulties_1_cm_nx511, 
         chipmulties_1_cm_nx513, chipmulties_1_cm_nx518, chipmulties_1_cm_nx523, 
         chipmulties_1_cm_nx528, chipmulties_1_cm_nx533, chipmulties_1_cm_nx535, 
         chipmulties_1_cm_nx537, chipmulties_1_cm_nx539, chipmulties_1_cm_nx541, 
         chipmulties_1_cm_nx543, chipmulties_1_cm_nx545, chipmulties_1_cm_nx547, 
         chipmulties_1_cm_nx550, chipmulties_1_cm_nx553, chipmulties_1_cm_nx555, 
         chipmulties_1_cm_nx557, chipmulties_1_cm_nx560, chipmulties_1_cm_nx562, 
         chipmulties_1_cm_nx566, chipmulties_1_cm_nx569, chipmulties_1_cm_nx571, 
         chipmulties_1_cm_nx573, chipmulties_1_cm_nx575, chipmulties_1_cm_nx580, 
         chipmulties_1_cm_nx583, chipmulties_1_cm_nx587, chipmulties_1_cm_nx589, 
         chipmulties_1_cm_nx591, chipmulties_0_cm_nx2, chipmulties_0_cm_nx10, 
         chipmulties_0_cm_nx12, chipmulties_0_cm_nx14, chipmulties_0_cm_nx18, 
         chipmulties_0_cm_nx22, chipmulties_0_cm_nx28, chipmulties_0_cm_nx46, 
         chipmulties_0_cm_nx52, chipmulties_0_cm_nx54, chipmulties_0_cm_nx62, 
         chipmulties_0_cm_nx68, chipmulties_0_cm_nx78, chipmulties_0_cm_nx118, 
         chipmulties_0_cm_nx130, chipmulties_0_cm_nx154, chipmulties_0_cm_nx164, 
         chipmulties_0_cm_nx178, chipmulties_0_cm_nx192, chipmulties_0_cm_nx228, 
         chipmulties_0_cm_nx501, chipmulties_0_cm_nx503, chipmulties_0_cm_nx506, 
         chipmulties_0_cm_nx508, chipmulties_0_cm_nx511, chipmulties_0_cm_nx513, 
         chipmulties_0_cm_nx518, chipmulties_0_cm_nx523, chipmulties_0_cm_nx528, 
         chipmulties_0_cm_nx533, chipmulties_0_cm_nx535, chipmulties_0_cm_nx537, 
         chipmulties_0_cm_nx539, chipmulties_0_cm_nx541, chipmulties_0_cm_nx543, 
         chipmulties_0_cm_nx545, chipmulties_0_cm_nx547, chipmulties_0_cm_nx550, 
         chipmulties_0_cm_nx553, chipmulties_0_cm_nx555, chipmulties_0_cm_nx557, 
         chipmulties_0_cm_nx560, chipmulties_0_cm_nx562, chipmulties_0_cm_nx566, 
         chipmulties_0_cm_nx569, chipmulties_0_cm_nx571, chipmulties_0_cm_nx573, 
         chipmulties_0_cm_nx575, chipmulties_0_cm_nx580, chipmulties_0_cm_nx583, 
         chipmulties_0_cm_nx587, chipmulties_0_cm_nx589, chipmulties_0_cm_nx591;



    nor04 chipmulties_15_cm_ix41 (.Y (C_15__0), .A0 (chipmulties_15_cm_nx501), .A1 (
          chipmulties_15_cm_nx503), .A2 (chipmulties_15_cm_nx508), .A3 (
          chipmulties_15_cm_nx518)) ;
    inv01 chipmulties_15_cm_ix502 (.Y (chipmulties_15_cm_nx501), .A (A_15__0)) ;
    oai21 chipmulties_15_cm_ix504 (.Y (chipmulties_15_cm_nx503), .A0 (
          chipmulties_15_cm_nx2), .A1 (A_15__2), .B0 (B_15__0)) ;
    nand02 chipmulties_15_cm_ix3 (.Y (chipmulties_15_cm_nx2), .A0 (
           chipmulties_15_cm_nx506), .A1 (A_15__4)) ;
    inv01 chipmulties_15_cm_ix507 (.Y (chipmulties_15_cm_nx506), .A (A_15__3)) ;
    oai21 chipmulties_15_cm_ix509 (.Y (chipmulties_15_cm_nx508), .A0 (
          chipmulties_15_cm_nx2), .A1 (A_15__1), .B0 (chipmulties_15_cm_nx28)) ;
    aoi21 chipmulties_15_cm_ix29 (.Y (chipmulties_15_cm_nx28), .A0 (
          chipmulties_15_cm_nx511), .A1 (A_15__2), .B0 (chipmulties_15_cm_nx513)
          ) ;
    nand03 chipmulties_15_cm_ix514 (.Y (chipmulties_15_cm_nx513), .A0 (
           chipmulties_15_cm_nx10), .A1 (chipmulties_15_cm_nx12), .A2 (
           chipmulties_15_cm_nx14)) ;
    xnor2 chipmulties_15_cm_ix11 (.Y (chipmulties_15_cm_nx10), .A0 (B_15__3), .A1 (
          B_15__4)) ;
    xnor2 chipmulties_15_cm_ix13 (.Y (chipmulties_15_cm_nx12), .A0 (B_15__2), .A1 (
          B_15__1)) ;
    xnor2 chipmulties_15_cm_ix15 (.Y (chipmulties_15_cm_nx14), .A0 (B_15__3), .A1 (
          B_15__2)) ;
    nor02 chipmulties_15_cm_ix75 (.Y (C_15__1), .A0 (chipmulties_15_cm_nx503), .A1 (
          chipmulties_15_cm_nx523)) ;
    aoi32 chipmulties_15_cm_ix524 (.Y (chipmulties_15_cm_nx523), .A0 (
          chipmulties_15_cm_nx52), .A1 (chipmulties_15_cm_nx54), .A2 (
          chipmulties_15_cm_nx28), .B0 (chipmulties_15_cm_nx46), .B1 (
          chipmulties_15_cm_nx68)) ;
    nor02 chipmulties_15_cm_ix53 (.Y (chipmulties_15_cm_nx52), .A0 (B_15__1), .A1 (
          chipmulties_15_cm_nx46)) ;
    nand02 chipmulties_15_cm_ix47 (.Y (chipmulties_15_cm_nx46), .A0 (A_15__0), .A1 (
           A_15__1)) ;
    nand02 chipmulties_15_cm_ix55 (.Y (chipmulties_15_cm_nx54), .A0 (
           chipmulties_15_cm_nx511), .A1 (chipmulties_15_cm_nx528)) ;
    inv01 chipmulties_15_cm_ix529 (.Y (chipmulties_15_cm_nx528), .A (B_15__4)) ;
    ao32 chipmulties_15_cm_ix69 (.Y (chipmulties_15_cm_nx68), .A0 (B_15__1), .A1 (
         A_15__0), .A2 (chipmulties_15_cm_nx62), .B0 (A_15__1), .B1 (
         chipmulties_15_cm_nx28)) ;
    aoi21 chipmulties_15_cm_ix63 (.Y (chipmulties_15_cm_nx62), .A0 (
          chipmulties_15_cm_nx511), .A1 (chipmulties_15_cm_nx528), .B0 (
          chipmulties_15_cm_nx508)) ;
    nor04 chipmulties_15_cm_ix109 (.Y (C_15__2), .A0 (chipmulties_15_cm_nx508), 
          .A1 (chipmulties_15_cm_nx533), .A2 (chipmulties_15_cm_nx535), .A3 (
          chipmulties_15_cm_nx537)) ;
    inv01 chipmulties_15_cm_ix534 (.Y (chipmulties_15_cm_nx533), .A (B_15__0)) ;
    nor03 chipmulties_15_cm_ix536 (.Y (chipmulties_15_cm_nx535), .A0 (A_15__0), 
          .A1 (A_15__1), .A2 (A_15__2)) ;
    ao22 chipmulties_15_cm_ix538 (.Y (chipmulties_15_cm_nx537), .A0 (
         chipmulties_15_cm_nx539), .A1 (chipmulties_15_cm_nx543), .B0 (
         chipmulties_15_cm_nx545), .B1 (chipmulties_15_cm_nx547)) ;
    oai21 chipmulties_15_cm_ix540 (.Y (chipmulties_15_cm_nx539), .A0 (A_15__2), 
          .A1 (B_15__1), .B0 (chipmulties_15_cm_nx541)) ;
    nor02 chipmulties_15_cm_ix542 (.Y (chipmulties_15_cm_nx541), .A0 (A_15__0), 
          .A1 (A_15__1)) ;
    xnor2 chipmulties_15_cm_ix544 (.Y (chipmulties_15_cm_nx543), .A0 (B_15__1), 
          .A1 (A_15__2)) ;
    oai22 chipmulties_15_cm_ix546 (.Y (chipmulties_15_cm_nx545), .A0 (
          chipmulties_15_cm_nx2), .A1 (chipmulties_15_cm_nx528), .B0 (
          chipmulties_15_cm_nx506), .B1 (A_15__4)) ;
    nand03 chipmulties_15_cm_ix548 (.Y (chipmulties_15_cm_nx547), .A0 (
           chipmulties_15_cm_nx2), .A1 (B_15__4), .A2 (chipmulties_15_cm_nx46)
           ) ;
    aoi21 chipmulties_15_cm_ix185 (.Y (C_15__3), .A0 (chipmulties_15_cm_nx550), 
          .A1 (chipmulties_15_cm_nx569), .B0 (chipmulties_15_cm_nx575)) ;
    oai21 chipmulties_15_cm_ix551 (.Y (chipmulties_15_cm_nx550), .A0 (
          chipmulties_15_cm_nx2), .A1 (A_15__1), .B0 (chipmulties_15_cm_nx178)
          ) ;
    oai22 chipmulties_15_cm_ix179 (.Y (chipmulties_15_cm_nx178), .A0 (
          chipmulties_15_cm_nx553), .A1 (chipmulties_15_cm_nx557), .B0 (
          chipmulties_15_cm_nx528), .B1 (chipmulties_15_cm_nx566)) ;
    aoi21 chipmulties_15_cm_ix554 (.Y (chipmulties_15_cm_nx553), .A0 (
          chipmulties_15_cm_nx555), .A1 (chipmulties_15_cm_nx46), .B0 (A_15__4)
          ) ;
    inv01 chipmulties_15_cm_ix556 (.Y (chipmulties_15_cm_nx555), .A (A_15__2)) ;
    nand02 chipmulties_15_cm_ix558 (.Y (chipmulties_15_cm_nx557), .A0 (
           chipmulties_15_cm_nx528), .A1 (chipmulties_15_cm_nx154)) ;
    oai21 chipmulties_15_cm_ix155 (.Y (chipmulties_15_cm_nx154), .A0 (
          chipmulties_15_cm_nx506), .A1 (A_15__0), .B0 (chipmulties_15_cm_nx560)
          ) ;
    aoi22 chipmulties_15_cm_ix561 (.Y (chipmulties_15_cm_nx560), .A0 (
          chipmulties_15_cm_nx562), .A1 (A_15__3), .B0 (chipmulties_15_cm_nx78)
          , .B1 (chipmulties_15_cm_nx130)) ;
    inv01 chipmulties_15_cm_ix563 (.Y (chipmulties_15_cm_nx562), .A (B_15__1)) ;
    aoi32 chipmulties_15_cm_ix567 (.Y (chipmulties_15_cm_nx566), .A0 (
          chipmulties_15_cm_nx164), .A1 (chipmulties_15_cm_nx78), .A2 (
          chipmulties_15_cm_nx130), .B0 (A_15__3), .B1 (chipmulties_15_cm_nx541)
          ) ;
    nand02 chipmulties_15_cm_ix165 (.Y (chipmulties_15_cm_nx164), .A0 (
           chipmulties_15_cm_nx555), .A1 (A_15__4)) ;
    or04 chipmulties_15_cm_ix570 (.Y (chipmulties_15_cm_nx569), .A0 (
         chipmulties_15_cm_nx528), .A1 (A_15__1), .A2 (chipmulties_15_cm_nx560)
         , .A3 (chipmulties_15_cm_nx571)) ;
    inv01 chipmulties_15_cm_ix574 (.Y (chipmulties_15_cm_nx573), .A (A_15__4)) ;
    nand03 chipmulties_15_cm_ix576 (.Y (chipmulties_15_cm_nx575), .A0 (
           chipmulties_15_cm_nx118), .A1 (B_15__0), .A2 (chipmulties_15_cm_nx18)
           ) ;
    nand03 chipmulties_15_cm_ix119 (.Y (chipmulties_15_cm_nx118), .A0 (B_15__4)
           , .A1 (A_15__2), .A2 (A_15__3)) ;
    nor02 chipmulties_15_cm_ix233 (.Y (C_15__4), .A0 (chipmulties_15_cm_nx575), 
          .A1 (chipmulties_15_cm_nx580)) ;
    aoi21 chipmulties_15_cm_ix581 (.Y (chipmulties_15_cm_nx580), .A0 (B_15__1), 
          .A1 (chipmulties_15_cm_nx192), .B0 (chipmulties_15_cm_nx228)) ;
    aoi21 chipmulties_15_cm_ix193 (.Y (chipmulties_15_cm_nx192), .A0 (
          chipmulties_15_cm_nx583), .A1 (B_15__4), .B0 (chipmulties_15_cm_nx22)
          ) ;
    oai33 chipmulties_15_cm_ix229 (.Y (chipmulties_15_cm_nx228), .A0 (
          chipmulties_15_cm_nx587), .A1 (chipmulties_15_cm_nx535), .A2 (
          chipmulties_15_cm_nx589), .B0 (B_15__1), .B1 (chipmulties_15_cm_nx573)
          , .B2 (chipmulties_15_cm_nx591)) ;
    aoi22 chipmulties_15_cm_ix588 (.Y (chipmulties_15_cm_nx587), .A0 (
          chipmulties_15_cm_nx562), .A1 (chipmulties_15_cm_nx571), .B0 (
          chipmulties_15_cm_nx573), .B1 (chipmulties_15_cm_nx130)) ;
    aoi21 chipmulties_15_cm_ix590 (.Y (chipmulties_15_cm_nx589), .A0 (A_15__2), 
          .A1 (A_15__1), .B0 (B_15__4)) ;
    oai21 chipmulties_15_cm_ix592 (.Y (chipmulties_15_cm_nx591), .A0 (
          chipmulties_15_cm_nx46), .A1 (chipmulties_15_cm_nx528), .B0 (A_15__3)
          ) ;
    inv01 chipmulties_15_cm_ix79 (.Y (chipmulties_15_cm_nx78), .A (
          chipmulties_15_cm_nx535)) ;
    inv01 chipmulties_15_cm_ix584 (.Y (chipmulties_15_cm_nx583), .A (
          chipmulties_15_cm_nx46)) ;
    inv01 chipmulties_15_cm_ix23 (.Y (chipmulties_15_cm_nx22), .A (
          chipmulties_15_cm_nx511)) ;
    inv01 chipmulties_15_cm_ix19 (.Y (chipmulties_15_cm_nx18), .A (
          chipmulties_15_cm_nx513)) ;
    inv01 chipmulties_15_cm_ix572 (.Y (chipmulties_15_cm_nx571), .A (
          chipmulties_15_cm_nx2)) ;
    nor02ii chipmulties_15_cm_ix512 (.Y (chipmulties_15_cm_nx511), .A0 (A_15__4)
            , .A1 (A_15__3)) ;
    and03 chipmulties_15_cm_ix519 (.Y (chipmulties_15_cm_nx518), .A0 (A_15__3), 
          .A1 (chipmulties_15_cm_nx573), .A2 (A_15__1)) ;
    nor02ii chipmulties_15_cm_ix131 (.Y (chipmulties_15_cm_nx130), .A0 (A_15__3)
            , .A1 (B_15__1)) ;
    nor04 chipmulties_14_cm_ix41 (.Y (C_14__0), .A0 (chipmulties_14_cm_nx501), .A1 (
          chipmulties_14_cm_nx503), .A2 (chipmulties_14_cm_nx508), .A3 (
          chipmulties_14_cm_nx518)) ;
    inv01 chipmulties_14_cm_ix502 (.Y (chipmulties_14_cm_nx501), .A (A_14__0)) ;
    oai21 chipmulties_14_cm_ix504 (.Y (chipmulties_14_cm_nx503), .A0 (
          chipmulties_14_cm_nx2), .A1 (A_14__2), .B0 (B_14__0)) ;
    nand02 chipmulties_14_cm_ix3 (.Y (chipmulties_14_cm_nx2), .A0 (
           chipmulties_14_cm_nx506), .A1 (A_14__4)) ;
    inv01 chipmulties_14_cm_ix507 (.Y (chipmulties_14_cm_nx506), .A (A_14__3)) ;
    oai21 chipmulties_14_cm_ix509 (.Y (chipmulties_14_cm_nx508), .A0 (
          chipmulties_14_cm_nx2), .A1 (A_14__1), .B0 (chipmulties_14_cm_nx28)) ;
    aoi21 chipmulties_14_cm_ix29 (.Y (chipmulties_14_cm_nx28), .A0 (
          chipmulties_14_cm_nx511), .A1 (A_14__2), .B0 (chipmulties_14_cm_nx513)
          ) ;
    nand03 chipmulties_14_cm_ix514 (.Y (chipmulties_14_cm_nx513), .A0 (
           chipmulties_14_cm_nx10), .A1 (chipmulties_14_cm_nx12), .A2 (
           chipmulties_14_cm_nx14)) ;
    xnor2 chipmulties_14_cm_ix11 (.Y (chipmulties_14_cm_nx10), .A0 (B_14__3), .A1 (
          B_14__4)) ;
    xnor2 chipmulties_14_cm_ix13 (.Y (chipmulties_14_cm_nx12), .A0 (B_14__2), .A1 (
          B_14__1)) ;
    xnor2 chipmulties_14_cm_ix15 (.Y (chipmulties_14_cm_nx14), .A0 (B_14__3), .A1 (
          B_14__2)) ;
    nor02 chipmulties_14_cm_ix75 (.Y (C_14__1), .A0 (chipmulties_14_cm_nx503), .A1 (
          chipmulties_14_cm_nx523)) ;
    aoi32 chipmulties_14_cm_ix524 (.Y (chipmulties_14_cm_nx523), .A0 (
          chipmulties_14_cm_nx52), .A1 (chipmulties_14_cm_nx54), .A2 (
          chipmulties_14_cm_nx28), .B0 (chipmulties_14_cm_nx46), .B1 (
          chipmulties_14_cm_nx68)) ;
    nor02 chipmulties_14_cm_ix53 (.Y (chipmulties_14_cm_nx52), .A0 (B_14__1), .A1 (
          chipmulties_14_cm_nx46)) ;
    nand02 chipmulties_14_cm_ix47 (.Y (chipmulties_14_cm_nx46), .A0 (A_14__0), .A1 (
           A_14__1)) ;
    nand02 chipmulties_14_cm_ix55 (.Y (chipmulties_14_cm_nx54), .A0 (
           chipmulties_14_cm_nx511), .A1 (chipmulties_14_cm_nx528)) ;
    inv01 chipmulties_14_cm_ix529 (.Y (chipmulties_14_cm_nx528), .A (B_14__4)) ;
    ao32 chipmulties_14_cm_ix69 (.Y (chipmulties_14_cm_nx68), .A0 (B_14__1), .A1 (
         A_14__0), .A2 (chipmulties_14_cm_nx62), .B0 (A_14__1), .B1 (
         chipmulties_14_cm_nx28)) ;
    aoi21 chipmulties_14_cm_ix63 (.Y (chipmulties_14_cm_nx62), .A0 (
          chipmulties_14_cm_nx511), .A1 (chipmulties_14_cm_nx528), .B0 (
          chipmulties_14_cm_nx508)) ;
    nor04 chipmulties_14_cm_ix109 (.Y (C_14__2), .A0 (chipmulties_14_cm_nx508), 
          .A1 (chipmulties_14_cm_nx533), .A2 (chipmulties_14_cm_nx535), .A3 (
          chipmulties_14_cm_nx537)) ;
    inv01 chipmulties_14_cm_ix534 (.Y (chipmulties_14_cm_nx533), .A (B_14__0)) ;
    nor03 chipmulties_14_cm_ix536 (.Y (chipmulties_14_cm_nx535), .A0 (A_14__0), 
          .A1 (A_14__1), .A2 (A_14__2)) ;
    ao22 chipmulties_14_cm_ix538 (.Y (chipmulties_14_cm_nx537), .A0 (
         chipmulties_14_cm_nx539), .A1 (chipmulties_14_cm_nx543), .B0 (
         chipmulties_14_cm_nx545), .B1 (chipmulties_14_cm_nx547)) ;
    oai21 chipmulties_14_cm_ix540 (.Y (chipmulties_14_cm_nx539), .A0 (A_14__2), 
          .A1 (B_14__1), .B0 (chipmulties_14_cm_nx541)) ;
    nor02 chipmulties_14_cm_ix542 (.Y (chipmulties_14_cm_nx541), .A0 (A_14__0), 
          .A1 (A_14__1)) ;
    xnor2 chipmulties_14_cm_ix544 (.Y (chipmulties_14_cm_nx543), .A0 (B_14__1), 
          .A1 (A_14__2)) ;
    oai22 chipmulties_14_cm_ix546 (.Y (chipmulties_14_cm_nx545), .A0 (
          chipmulties_14_cm_nx2), .A1 (chipmulties_14_cm_nx528), .B0 (
          chipmulties_14_cm_nx506), .B1 (A_14__4)) ;
    nand03 chipmulties_14_cm_ix548 (.Y (chipmulties_14_cm_nx547), .A0 (
           chipmulties_14_cm_nx2), .A1 (B_14__4), .A2 (chipmulties_14_cm_nx46)
           ) ;
    aoi21 chipmulties_14_cm_ix185 (.Y (C_14__3), .A0 (chipmulties_14_cm_nx550), 
          .A1 (chipmulties_14_cm_nx569), .B0 (chipmulties_14_cm_nx575)) ;
    oai21 chipmulties_14_cm_ix551 (.Y (chipmulties_14_cm_nx550), .A0 (
          chipmulties_14_cm_nx2), .A1 (A_14__1), .B0 (chipmulties_14_cm_nx178)
          ) ;
    oai22 chipmulties_14_cm_ix179 (.Y (chipmulties_14_cm_nx178), .A0 (
          chipmulties_14_cm_nx553), .A1 (chipmulties_14_cm_nx557), .B0 (
          chipmulties_14_cm_nx528), .B1 (chipmulties_14_cm_nx566)) ;
    aoi21 chipmulties_14_cm_ix554 (.Y (chipmulties_14_cm_nx553), .A0 (
          chipmulties_14_cm_nx555), .A1 (chipmulties_14_cm_nx46), .B0 (A_14__4)
          ) ;
    inv01 chipmulties_14_cm_ix556 (.Y (chipmulties_14_cm_nx555), .A (A_14__2)) ;
    nand02 chipmulties_14_cm_ix558 (.Y (chipmulties_14_cm_nx557), .A0 (
           chipmulties_14_cm_nx528), .A1 (chipmulties_14_cm_nx154)) ;
    oai21 chipmulties_14_cm_ix155 (.Y (chipmulties_14_cm_nx154), .A0 (
          chipmulties_14_cm_nx506), .A1 (A_14__0), .B0 (chipmulties_14_cm_nx560)
          ) ;
    aoi22 chipmulties_14_cm_ix561 (.Y (chipmulties_14_cm_nx560), .A0 (
          chipmulties_14_cm_nx562), .A1 (A_14__3), .B0 (chipmulties_14_cm_nx78)
          , .B1 (chipmulties_14_cm_nx130)) ;
    inv01 chipmulties_14_cm_ix563 (.Y (chipmulties_14_cm_nx562), .A (B_14__1)) ;
    aoi32 chipmulties_14_cm_ix567 (.Y (chipmulties_14_cm_nx566), .A0 (
          chipmulties_14_cm_nx164), .A1 (chipmulties_14_cm_nx78), .A2 (
          chipmulties_14_cm_nx130), .B0 (A_14__3), .B1 (chipmulties_14_cm_nx541)
          ) ;
    nand02 chipmulties_14_cm_ix165 (.Y (chipmulties_14_cm_nx164), .A0 (
           chipmulties_14_cm_nx555), .A1 (A_14__4)) ;
    or04 chipmulties_14_cm_ix570 (.Y (chipmulties_14_cm_nx569), .A0 (
         chipmulties_14_cm_nx528), .A1 (A_14__1), .A2 (chipmulties_14_cm_nx560)
         , .A3 (chipmulties_14_cm_nx571)) ;
    inv01 chipmulties_14_cm_ix574 (.Y (chipmulties_14_cm_nx573), .A (A_14__4)) ;
    nand03 chipmulties_14_cm_ix576 (.Y (chipmulties_14_cm_nx575), .A0 (
           chipmulties_14_cm_nx118), .A1 (B_14__0), .A2 (chipmulties_14_cm_nx18)
           ) ;
    nand03 chipmulties_14_cm_ix119 (.Y (chipmulties_14_cm_nx118), .A0 (B_14__4)
           , .A1 (A_14__2), .A2 (A_14__3)) ;
    nor02 chipmulties_14_cm_ix233 (.Y (C_14__4), .A0 (chipmulties_14_cm_nx575), 
          .A1 (chipmulties_14_cm_nx580)) ;
    aoi21 chipmulties_14_cm_ix581 (.Y (chipmulties_14_cm_nx580), .A0 (B_14__1), 
          .A1 (chipmulties_14_cm_nx192), .B0 (chipmulties_14_cm_nx228)) ;
    aoi21 chipmulties_14_cm_ix193 (.Y (chipmulties_14_cm_nx192), .A0 (
          chipmulties_14_cm_nx583), .A1 (B_14__4), .B0 (chipmulties_14_cm_nx22)
          ) ;
    oai33 chipmulties_14_cm_ix229 (.Y (chipmulties_14_cm_nx228), .A0 (
          chipmulties_14_cm_nx587), .A1 (chipmulties_14_cm_nx535), .A2 (
          chipmulties_14_cm_nx589), .B0 (B_14__1), .B1 (chipmulties_14_cm_nx573)
          , .B2 (chipmulties_14_cm_nx591)) ;
    aoi22 chipmulties_14_cm_ix588 (.Y (chipmulties_14_cm_nx587), .A0 (
          chipmulties_14_cm_nx562), .A1 (chipmulties_14_cm_nx571), .B0 (
          chipmulties_14_cm_nx573), .B1 (chipmulties_14_cm_nx130)) ;
    aoi21 chipmulties_14_cm_ix590 (.Y (chipmulties_14_cm_nx589), .A0 (A_14__2), 
          .A1 (A_14__1), .B0 (B_14__4)) ;
    oai21 chipmulties_14_cm_ix592 (.Y (chipmulties_14_cm_nx591), .A0 (
          chipmulties_14_cm_nx46), .A1 (chipmulties_14_cm_nx528), .B0 (A_14__3)
          ) ;
    inv01 chipmulties_14_cm_ix79 (.Y (chipmulties_14_cm_nx78), .A (
          chipmulties_14_cm_nx535)) ;
    inv01 chipmulties_14_cm_ix584 (.Y (chipmulties_14_cm_nx583), .A (
          chipmulties_14_cm_nx46)) ;
    inv01 chipmulties_14_cm_ix23 (.Y (chipmulties_14_cm_nx22), .A (
          chipmulties_14_cm_nx511)) ;
    inv01 chipmulties_14_cm_ix19 (.Y (chipmulties_14_cm_nx18), .A (
          chipmulties_14_cm_nx513)) ;
    inv01 chipmulties_14_cm_ix572 (.Y (chipmulties_14_cm_nx571), .A (
          chipmulties_14_cm_nx2)) ;
    nor02ii chipmulties_14_cm_ix512 (.Y (chipmulties_14_cm_nx511), .A0 (A_14__4)
            , .A1 (A_14__3)) ;
    and03 chipmulties_14_cm_ix519 (.Y (chipmulties_14_cm_nx518), .A0 (A_14__3), 
          .A1 (chipmulties_14_cm_nx573), .A2 (A_14__1)) ;
    nor02ii chipmulties_14_cm_ix131 (.Y (chipmulties_14_cm_nx130), .A0 (A_14__3)
            , .A1 (B_14__1)) ;
    nor04 chipmulties_13_cm_ix41 (.Y (C_13__0), .A0 (chipmulties_13_cm_nx501), .A1 (
          chipmulties_13_cm_nx503), .A2 (chipmulties_13_cm_nx508), .A3 (
          chipmulties_13_cm_nx518)) ;
    inv01 chipmulties_13_cm_ix502 (.Y (chipmulties_13_cm_nx501), .A (A_13__0)) ;
    oai21 chipmulties_13_cm_ix504 (.Y (chipmulties_13_cm_nx503), .A0 (
          chipmulties_13_cm_nx2), .A1 (A_13__2), .B0 (B_13__0)) ;
    nand02 chipmulties_13_cm_ix3 (.Y (chipmulties_13_cm_nx2), .A0 (
           chipmulties_13_cm_nx506), .A1 (A_13__4)) ;
    inv01 chipmulties_13_cm_ix507 (.Y (chipmulties_13_cm_nx506), .A (A_13__3)) ;
    oai21 chipmulties_13_cm_ix509 (.Y (chipmulties_13_cm_nx508), .A0 (
          chipmulties_13_cm_nx2), .A1 (A_13__1), .B0 (chipmulties_13_cm_nx28)) ;
    aoi21 chipmulties_13_cm_ix29 (.Y (chipmulties_13_cm_nx28), .A0 (
          chipmulties_13_cm_nx511), .A1 (A_13__2), .B0 (chipmulties_13_cm_nx513)
          ) ;
    nand03 chipmulties_13_cm_ix514 (.Y (chipmulties_13_cm_nx513), .A0 (
           chipmulties_13_cm_nx10), .A1 (chipmulties_13_cm_nx12), .A2 (
           chipmulties_13_cm_nx14)) ;
    xnor2 chipmulties_13_cm_ix11 (.Y (chipmulties_13_cm_nx10), .A0 (B_13__3), .A1 (
          B_13__4)) ;
    xnor2 chipmulties_13_cm_ix13 (.Y (chipmulties_13_cm_nx12), .A0 (B_13__2), .A1 (
          B_13__1)) ;
    xnor2 chipmulties_13_cm_ix15 (.Y (chipmulties_13_cm_nx14), .A0 (B_13__3), .A1 (
          B_13__2)) ;
    nor02 chipmulties_13_cm_ix75 (.Y (C_13__1), .A0 (chipmulties_13_cm_nx503), .A1 (
          chipmulties_13_cm_nx523)) ;
    aoi32 chipmulties_13_cm_ix524 (.Y (chipmulties_13_cm_nx523), .A0 (
          chipmulties_13_cm_nx52), .A1 (chipmulties_13_cm_nx54), .A2 (
          chipmulties_13_cm_nx28), .B0 (chipmulties_13_cm_nx46), .B1 (
          chipmulties_13_cm_nx68)) ;
    nor02 chipmulties_13_cm_ix53 (.Y (chipmulties_13_cm_nx52), .A0 (B_13__1), .A1 (
          chipmulties_13_cm_nx46)) ;
    nand02 chipmulties_13_cm_ix47 (.Y (chipmulties_13_cm_nx46), .A0 (A_13__0), .A1 (
           A_13__1)) ;
    nand02 chipmulties_13_cm_ix55 (.Y (chipmulties_13_cm_nx54), .A0 (
           chipmulties_13_cm_nx511), .A1 (chipmulties_13_cm_nx528)) ;
    inv01 chipmulties_13_cm_ix529 (.Y (chipmulties_13_cm_nx528), .A (B_13__4)) ;
    ao32 chipmulties_13_cm_ix69 (.Y (chipmulties_13_cm_nx68), .A0 (B_13__1), .A1 (
         A_13__0), .A2 (chipmulties_13_cm_nx62), .B0 (A_13__1), .B1 (
         chipmulties_13_cm_nx28)) ;
    aoi21 chipmulties_13_cm_ix63 (.Y (chipmulties_13_cm_nx62), .A0 (
          chipmulties_13_cm_nx511), .A1 (chipmulties_13_cm_nx528), .B0 (
          chipmulties_13_cm_nx508)) ;
    nor04 chipmulties_13_cm_ix109 (.Y (C_13__2), .A0 (chipmulties_13_cm_nx508), 
          .A1 (chipmulties_13_cm_nx533), .A2 (chipmulties_13_cm_nx535), .A3 (
          chipmulties_13_cm_nx537)) ;
    inv01 chipmulties_13_cm_ix534 (.Y (chipmulties_13_cm_nx533), .A (B_13__0)) ;
    nor03 chipmulties_13_cm_ix536 (.Y (chipmulties_13_cm_nx535), .A0 (A_13__0), 
          .A1 (A_13__1), .A2 (A_13__2)) ;
    ao22 chipmulties_13_cm_ix538 (.Y (chipmulties_13_cm_nx537), .A0 (
         chipmulties_13_cm_nx539), .A1 (chipmulties_13_cm_nx543), .B0 (
         chipmulties_13_cm_nx545), .B1 (chipmulties_13_cm_nx547)) ;
    oai21 chipmulties_13_cm_ix540 (.Y (chipmulties_13_cm_nx539), .A0 (A_13__2), 
          .A1 (B_13__1), .B0 (chipmulties_13_cm_nx541)) ;
    nor02 chipmulties_13_cm_ix542 (.Y (chipmulties_13_cm_nx541), .A0 (A_13__0), 
          .A1 (A_13__1)) ;
    xnor2 chipmulties_13_cm_ix544 (.Y (chipmulties_13_cm_nx543), .A0 (B_13__1), 
          .A1 (A_13__2)) ;
    oai22 chipmulties_13_cm_ix546 (.Y (chipmulties_13_cm_nx545), .A0 (
          chipmulties_13_cm_nx2), .A1 (chipmulties_13_cm_nx528), .B0 (
          chipmulties_13_cm_nx506), .B1 (A_13__4)) ;
    nand03 chipmulties_13_cm_ix548 (.Y (chipmulties_13_cm_nx547), .A0 (
           chipmulties_13_cm_nx2), .A1 (B_13__4), .A2 (chipmulties_13_cm_nx46)
           ) ;
    aoi21 chipmulties_13_cm_ix185 (.Y (C_13__3), .A0 (chipmulties_13_cm_nx550), 
          .A1 (chipmulties_13_cm_nx569), .B0 (chipmulties_13_cm_nx575)) ;
    oai21 chipmulties_13_cm_ix551 (.Y (chipmulties_13_cm_nx550), .A0 (
          chipmulties_13_cm_nx2), .A1 (A_13__1), .B0 (chipmulties_13_cm_nx178)
          ) ;
    oai22 chipmulties_13_cm_ix179 (.Y (chipmulties_13_cm_nx178), .A0 (
          chipmulties_13_cm_nx553), .A1 (chipmulties_13_cm_nx557), .B0 (
          chipmulties_13_cm_nx528), .B1 (chipmulties_13_cm_nx566)) ;
    aoi21 chipmulties_13_cm_ix554 (.Y (chipmulties_13_cm_nx553), .A0 (
          chipmulties_13_cm_nx555), .A1 (chipmulties_13_cm_nx46), .B0 (A_13__4)
          ) ;
    inv01 chipmulties_13_cm_ix556 (.Y (chipmulties_13_cm_nx555), .A (A_13__2)) ;
    nand02 chipmulties_13_cm_ix558 (.Y (chipmulties_13_cm_nx557), .A0 (
           chipmulties_13_cm_nx528), .A1 (chipmulties_13_cm_nx154)) ;
    oai21 chipmulties_13_cm_ix155 (.Y (chipmulties_13_cm_nx154), .A0 (
          chipmulties_13_cm_nx506), .A1 (A_13__0), .B0 (chipmulties_13_cm_nx560)
          ) ;
    aoi22 chipmulties_13_cm_ix561 (.Y (chipmulties_13_cm_nx560), .A0 (
          chipmulties_13_cm_nx562), .A1 (A_13__3), .B0 (chipmulties_13_cm_nx78)
          , .B1 (chipmulties_13_cm_nx130)) ;
    inv01 chipmulties_13_cm_ix563 (.Y (chipmulties_13_cm_nx562), .A (B_13__1)) ;
    aoi32 chipmulties_13_cm_ix567 (.Y (chipmulties_13_cm_nx566), .A0 (
          chipmulties_13_cm_nx164), .A1 (chipmulties_13_cm_nx78), .A2 (
          chipmulties_13_cm_nx130), .B0 (A_13__3), .B1 (chipmulties_13_cm_nx541)
          ) ;
    nand02 chipmulties_13_cm_ix165 (.Y (chipmulties_13_cm_nx164), .A0 (
           chipmulties_13_cm_nx555), .A1 (A_13__4)) ;
    or04 chipmulties_13_cm_ix570 (.Y (chipmulties_13_cm_nx569), .A0 (
         chipmulties_13_cm_nx528), .A1 (A_13__1), .A2 (chipmulties_13_cm_nx560)
         , .A3 (chipmulties_13_cm_nx571)) ;
    inv01 chipmulties_13_cm_ix574 (.Y (chipmulties_13_cm_nx573), .A (A_13__4)) ;
    nand03 chipmulties_13_cm_ix576 (.Y (chipmulties_13_cm_nx575), .A0 (
           chipmulties_13_cm_nx118), .A1 (B_13__0), .A2 (chipmulties_13_cm_nx18)
           ) ;
    nand03 chipmulties_13_cm_ix119 (.Y (chipmulties_13_cm_nx118), .A0 (B_13__4)
           , .A1 (A_13__2), .A2 (A_13__3)) ;
    nor02 chipmulties_13_cm_ix233 (.Y (C_13__4), .A0 (chipmulties_13_cm_nx575), 
          .A1 (chipmulties_13_cm_nx580)) ;
    aoi21 chipmulties_13_cm_ix581 (.Y (chipmulties_13_cm_nx580), .A0 (B_13__1), 
          .A1 (chipmulties_13_cm_nx192), .B0 (chipmulties_13_cm_nx228)) ;
    aoi21 chipmulties_13_cm_ix193 (.Y (chipmulties_13_cm_nx192), .A0 (
          chipmulties_13_cm_nx583), .A1 (B_13__4), .B0 (chipmulties_13_cm_nx22)
          ) ;
    oai33 chipmulties_13_cm_ix229 (.Y (chipmulties_13_cm_nx228), .A0 (
          chipmulties_13_cm_nx587), .A1 (chipmulties_13_cm_nx535), .A2 (
          chipmulties_13_cm_nx589), .B0 (B_13__1), .B1 (chipmulties_13_cm_nx573)
          , .B2 (chipmulties_13_cm_nx591)) ;
    aoi22 chipmulties_13_cm_ix588 (.Y (chipmulties_13_cm_nx587), .A0 (
          chipmulties_13_cm_nx562), .A1 (chipmulties_13_cm_nx571), .B0 (
          chipmulties_13_cm_nx573), .B1 (chipmulties_13_cm_nx130)) ;
    aoi21 chipmulties_13_cm_ix590 (.Y (chipmulties_13_cm_nx589), .A0 (A_13__2), 
          .A1 (A_13__1), .B0 (B_13__4)) ;
    oai21 chipmulties_13_cm_ix592 (.Y (chipmulties_13_cm_nx591), .A0 (
          chipmulties_13_cm_nx46), .A1 (chipmulties_13_cm_nx528), .B0 (A_13__3)
          ) ;
    inv01 chipmulties_13_cm_ix79 (.Y (chipmulties_13_cm_nx78), .A (
          chipmulties_13_cm_nx535)) ;
    inv01 chipmulties_13_cm_ix584 (.Y (chipmulties_13_cm_nx583), .A (
          chipmulties_13_cm_nx46)) ;
    inv01 chipmulties_13_cm_ix23 (.Y (chipmulties_13_cm_nx22), .A (
          chipmulties_13_cm_nx511)) ;
    inv01 chipmulties_13_cm_ix19 (.Y (chipmulties_13_cm_nx18), .A (
          chipmulties_13_cm_nx513)) ;
    inv01 chipmulties_13_cm_ix572 (.Y (chipmulties_13_cm_nx571), .A (
          chipmulties_13_cm_nx2)) ;
    nor02ii chipmulties_13_cm_ix512 (.Y (chipmulties_13_cm_nx511), .A0 (A_13__4)
            , .A1 (A_13__3)) ;
    and03 chipmulties_13_cm_ix519 (.Y (chipmulties_13_cm_nx518), .A0 (A_13__3), 
          .A1 (chipmulties_13_cm_nx573), .A2 (A_13__1)) ;
    nor02ii chipmulties_13_cm_ix131 (.Y (chipmulties_13_cm_nx130), .A0 (A_13__3)
            , .A1 (B_13__1)) ;
    nor04 chipmulties_12_cm_ix41 (.Y (C_12__0), .A0 (chipmulties_12_cm_nx501), .A1 (
          chipmulties_12_cm_nx503), .A2 (chipmulties_12_cm_nx508), .A3 (
          chipmulties_12_cm_nx518)) ;
    inv01 chipmulties_12_cm_ix502 (.Y (chipmulties_12_cm_nx501), .A (A_12__0)) ;
    oai21 chipmulties_12_cm_ix504 (.Y (chipmulties_12_cm_nx503), .A0 (
          chipmulties_12_cm_nx2), .A1 (A_12__2), .B0 (B_12__0)) ;
    nand02 chipmulties_12_cm_ix3 (.Y (chipmulties_12_cm_nx2), .A0 (
           chipmulties_12_cm_nx506), .A1 (A_12__4)) ;
    inv01 chipmulties_12_cm_ix507 (.Y (chipmulties_12_cm_nx506), .A (A_12__3)) ;
    oai21 chipmulties_12_cm_ix509 (.Y (chipmulties_12_cm_nx508), .A0 (
          chipmulties_12_cm_nx2), .A1 (A_12__1), .B0 (chipmulties_12_cm_nx28)) ;
    aoi21 chipmulties_12_cm_ix29 (.Y (chipmulties_12_cm_nx28), .A0 (
          chipmulties_12_cm_nx511), .A1 (A_12__2), .B0 (chipmulties_12_cm_nx513)
          ) ;
    nand03 chipmulties_12_cm_ix514 (.Y (chipmulties_12_cm_nx513), .A0 (
           chipmulties_12_cm_nx10), .A1 (chipmulties_12_cm_nx12), .A2 (
           chipmulties_12_cm_nx14)) ;
    xnor2 chipmulties_12_cm_ix11 (.Y (chipmulties_12_cm_nx10), .A0 (B_12__3), .A1 (
          B_12__4)) ;
    xnor2 chipmulties_12_cm_ix13 (.Y (chipmulties_12_cm_nx12), .A0 (B_12__2), .A1 (
          B_12__1)) ;
    xnor2 chipmulties_12_cm_ix15 (.Y (chipmulties_12_cm_nx14), .A0 (B_12__3), .A1 (
          B_12__2)) ;
    nor02 chipmulties_12_cm_ix75 (.Y (C_12__1), .A0 (chipmulties_12_cm_nx503), .A1 (
          chipmulties_12_cm_nx523)) ;
    aoi32 chipmulties_12_cm_ix524 (.Y (chipmulties_12_cm_nx523), .A0 (
          chipmulties_12_cm_nx52), .A1 (chipmulties_12_cm_nx54), .A2 (
          chipmulties_12_cm_nx28), .B0 (chipmulties_12_cm_nx46), .B1 (
          chipmulties_12_cm_nx68)) ;
    nor02 chipmulties_12_cm_ix53 (.Y (chipmulties_12_cm_nx52), .A0 (B_12__1), .A1 (
          chipmulties_12_cm_nx46)) ;
    nand02 chipmulties_12_cm_ix47 (.Y (chipmulties_12_cm_nx46), .A0 (A_12__0), .A1 (
           A_12__1)) ;
    nand02 chipmulties_12_cm_ix55 (.Y (chipmulties_12_cm_nx54), .A0 (
           chipmulties_12_cm_nx511), .A1 (chipmulties_12_cm_nx528)) ;
    inv01 chipmulties_12_cm_ix529 (.Y (chipmulties_12_cm_nx528), .A (B_12__4)) ;
    ao32 chipmulties_12_cm_ix69 (.Y (chipmulties_12_cm_nx68), .A0 (B_12__1), .A1 (
         A_12__0), .A2 (chipmulties_12_cm_nx62), .B0 (A_12__1), .B1 (
         chipmulties_12_cm_nx28)) ;
    aoi21 chipmulties_12_cm_ix63 (.Y (chipmulties_12_cm_nx62), .A0 (
          chipmulties_12_cm_nx511), .A1 (chipmulties_12_cm_nx528), .B0 (
          chipmulties_12_cm_nx508)) ;
    nor04 chipmulties_12_cm_ix109 (.Y (C_12__2), .A0 (chipmulties_12_cm_nx508), 
          .A1 (chipmulties_12_cm_nx533), .A2 (chipmulties_12_cm_nx535), .A3 (
          chipmulties_12_cm_nx537)) ;
    inv01 chipmulties_12_cm_ix534 (.Y (chipmulties_12_cm_nx533), .A (B_12__0)) ;
    nor03 chipmulties_12_cm_ix536 (.Y (chipmulties_12_cm_nx535), .A0 (A_12__0), 
          .A1 (A_12__1), .A2 (A_12__2)) ;
    ao22 chipmulties_12_cm_ix538 (.Y (chipmulties_12_cm_nx537), .A0 (
         chipmulties_12_cm_nx539), .A1 (chipmulties_12_cm_nx543), .B0 (
         chipmulties_12_cm_nx545), .B1 (chipmulties_12_cm_nx547)) ;
    oai21 chipmulties_12_cm_ix540 (.Y (chipmulties_12_cm_nx539), .A0 (A_12__2), 
          .A1 (B_12__1), .B0 (chipmulties_12_cm_nx541)) ;
    nor02 chipmulties_12_cm_ix542 (.Y (chipmulties_12_cm_nx541), .A0 (A_12__0), 
          .A1 (A_12__1)) ;
    xnor2 chipmulties_12_cm_ix544 (.Y (chipmulties_12_cm_nx543), .A0 (B_12__1), 
          .A1 (A_12__2)) ;
    oai22 chipmulties_12_cm_ix546 (.Y (chipmulties_12_cm_nx545), .A0 (
          chipmulties_12_cm_nx2), .A1 (chipmulties_12_cm_nx528), .B0 (
          chipmulties_12_cm_nx506), .B1 (A_12__4)) ;
    nand03 chipmulties_12_cm_ix548 (.Y (chipmulties_12_cm_nx547), .A0 (
           chipmulties_12_cm_nx2), .A1 (B_12__4), .A2 (chipmulties_12_cm_nx46)
           ) ;
    aoi21 chipmulties_12_cm_ix185 (.Y (C_12__3), .A0 (chipmulties_12_cm_nx550), 
          .A1 (chipmulties_12_cm_nx569), .B0 (chipmulties_12_cm_nx575)) ;
    oai21 chipmulties_12_cm_ix551 (.Y (chipmulties_12_cm_nx550), .A0 (
          chipmulties_12_cm_nx2), .A1 (A_12__1), .B0 (chipmulties_12_cm_nx178)
          ) ;
    oai22 chipmulties_12_cm_ix179 (.Y (chipmulties_12_cm_nx178), .A0 (
          chipmulties_12_cm_nx553), .A1 (chipmulties_12_cm_nx557), .B0 (
          chipmulties_12_cm_nx528), .B1 (chipmulties_12_cm_nx566)) ;
    aoi21 chipmulties_12_cm_ix554 (.Y (chipmulties_12_cm_nx553), .A0 (
          chipmulties_12_cm_nx555), .A1 (chipmulties_12_cm_nx46), .B0 (A_12__4)
          ) ;
    inv01 chipmulties_12_cm_ix556 (.Y (chipmulties_12_cm_nx555), .A (A_12__2)) ;
    nand02 chipmulties_12_cm_ix558 (.Y (chipmulties_12_cm_nx557), .A0 (
           chipmulties_12_cm_nx528), .A1 (chipmulties_12_cm_nx154)) ;
    oai21 chipmulties_12_cm_ix155 (.Y (chipmulties_12_cm_nx154), .A0 (
          chipmulties_12_cm_nx506), .A1 (A_12__0), .B0 (chipmulties_12_cm_nx560)
          ) ;
    aoi22 chipmulties_12_cm_ix561 (.Y (chipmulties_12_cm_nx560), .A0 (
          chipmulties_12_cm_nx562), .A1 (A_12__3), .B0 (chipmulties_12_cm_nx78)
          , .B1 (chipmulties_12_cm_nx130)) ;
    inv01 chipmulties_12_cm_ix563 (.Y (chipmulties_12_cm_nx562), .A (B_12__1)) ;
    aoi32 chipmulties_12_cm_ix567 (.Y (chipmulties_12_cm_nx566), .A0 (
          chipmulties_12_cm_nx164), .A1 (chipmulties_12_cm_nx78), .A2 (
          chipmulties_12_cm_nx130), .B0 (A_12__3), .B1 (chipmulties_12_cm_nx541)
          ) ;
    nand02 chipmulties_12_cm_ix165 (.Y (chipmulties_12_cm_nx164), .A0 (
           chipmulties_12_cm_nx555), .A1 (A_12__4)) ;
    or04 chipmulties_12_cm_ix570 (.Y (chipmulties_12_cm_nx569), .A0 (
         chipmulties_12_cm_nx528), .A1 (A_12__1), .A2 (chipmulties_12_cm_nx560)
         , .A3 (chipmulties_12_cm_nx571)) ;
    inv01 chipmulties_12_cm_ix574 (.Y (chipmulties_12_cm_nx573), .A (A_12__4)) ;
    nand03 chipmulties_12_cm_ix576 (.Y (chipmulties_12_cm_nx575), .A0 (
           chipmulties_12_cm_nx118), .A1 (B_12__0), .A2 (chipmulties_12_cm_nx18)
           ) ;
    nand03 chipmulties_12_cm_ix119 (.Y (chipmulties_12_cm_nx118), .A0 (B_12__4)
           , .A1 (A_12__2), .A2 (A_12__3)) ;
    nor02 chipmulties_12_cm_ix233 (.Y (C_12__4), .A0 (chipmulties_12_cm_nx575), 
          .A1 (chipmulties_12_cm_nx580)) ;
    aoi21 chipmulties_12_cm_ix581 (.Y (chipmulties_12_cm_nx580), .A0 (B_12__1), 
          .A1 (chipmulties_12_cm_nx192), .B0 (chipmulties_12_cm_nx228)) ;
    aoi21 chipmulties_12_cm_ix193 (.Y (chipmulties_12_cm_nx192), .A0 (
          chipmulties_12_cm_nx583), .A1 (B_12__4), .B0 (chipmulties_12_cm_nx22)
          ) ;
    oai33 chipmulties_12_cm_ix229 (.Y (chipmulties_12_cm_nx228), .A0 (
          chipmulties_12_cm_nx587), .A1 (chipmulties_12_cm_nx535), .A2 (
          chipmulties_12_cm_nx589), .B0 (B_12__1), .B1 (chipmulties_12_cm_nx573)
          , .B2 (chipmulties_12_cm_nx591)) ;
    aoi22 chipmulties_12_cm_ix588 (.Y (chipmulties_12_cm_nx587), .A0 (
          chipmulties_12_cm_nx562), .A1 (chipmulties_12_cm_nx571), .B0 (
          chipmulties_12_cm_nx573), .B1 (chipmulties_12_cm_nx130)) ;
    aoi21 chipmulties_12_cm_ix590 (.Y (chipmulties_12_cm_nx589), .A0 (A_12__2), 
          .A1 (A_12__1), .B0 (B_12__4)) ;
    oai21 chipmulties_12_cm_ix592 (.Y (chipmulties_12_cm_nx591), .A0 (
          chipmulties_12_cm_nx46), .A1 (chipmulties_12_cm_nx528), .B0 (A_12__3)
          ) ;
    inv01 chipmulties_12_cm_ix79 (.Y (chipmulties_12_cm_nx78), .A (
          chipmulties_12_cm_nx535)) ;
    inv01 chipmulties_12_cm_ix584 (.Y (chipmulties_12_cm_nx583), .A (
          chipmulties_12_cm_nx46)) ;
    inv01 chipmulties_12_cm_ix23 (.Y (chipmulties_12_cm_nx22), .A (
          chipmulties_12_cm_nx511)) ;
    inv01 chipmulties_12_cm_ix19 (.Y (chipmulties_12_cm_nx18), .A (
          chipmulties_12_cm_nx513)) ;
    inv01 chipmulties_12_cm_ix572 (.Y (chipmulties_12_cm_nx571), .A (
          chipmulties_12_cm_nx2)) ;
    nor02ii chipmulties_12_cm_ix512 (.Y (chipmulties_12_cm_nx511), .A0 (A_12__4)
            , .A1 (A_12__3)) ;
    and03 chipmulties_12_cm_ix519 (.Y (chipmulties_12_cm_nx518), .A0 (A_12__3), 
          .A1 (chipmulties_12_cm_nx573), .A2 (A_12__1)) ;
    nor02ii chipmulties_12_cm_ix131 (.Y (chipmulties_12_cm_nx130), .A0 (A_12__3)
            , .A1 (B_12__1)) ;
    nor04 chipmulties_11_cm_ix41 (.Y (C_11__0), .A0 (chipmulties_11_cm_nx501), .A1 (
          chipmulties_11_cm_nx503), .A2 (chipmulties_11_cm_nx508), .A3 (
          chipmulties_11_cm_nx518)) ;
    inv01 chipmulties_11_cm_ix502 (.Y (chipmulties_11_cm_nx501), .A (A_11__0)) ;
    oai21 chipmulties_11_cm_ix504 (.Y (chipmulties_11_cm_nx503), .A0 (
          chipmulties_11_cm_nx2), .A1 (A_11__2), .B0 (B_11__0)) ;
    nand02 chipmulties_11_cm_ix3 (.Y (chipmulties_11_cm_nx2), .A0 (
           chipmulties_11_cm_nx506), .A1 (A_11__4)) ;
    inv01 chipmulties_11_cm_ix507 (.Y (chipmulties_11_cm_nx506), .A (A_11__3)) ;
    oai21 chipmulties_11_cm_ix509 (.Y (chipmulties_11_cm_nx508), .A0 (
          chipmulties_11_cm_nx2), .A1 (A_11__1), .B0 (chipmulties_11_cm_nx28)) ;
    aoi21 chipmulties_11_cm_ix29 (.Y (chipmulties_11_cm_nx28), .A0 (
          chipmulties_11_cm_nx511), .A1 (A_11__2), .B0 (chipmulties_11_cm_nx513)
          ) ;
    nand03 chipmulties_11_cm_ix514 (.Y (chipmulties_11_cm_nx513), .A0 (
           chipmulties_11_cm_nx10), .A1 (chipmulties_11_cm_nx12), .A2 (
           chipmulties_11_cm_nx14)) ;
    xnor2 chipmulties_11_cm_ix11 (.Y (chipmulties_11_cm_nx10), .A0 (B_11__3), .A1 (
          B_11__4)) ;
    xnor2 chipmulties_11_cm_ix13 (.Y (chipmulties_11_cm_nx12), .A0 (B_11__2), .A1 (
          B_11__1)) ;
    xnor2 chipmulties_11_cm_ix15 (.Y (chipmulties_11_cm_nx14), .A0 (B_11__3), .A1 (
          B_11__2)) ;
    nor02 chipmulties_11_cm_ix75 (.Y (C_11__1), .A0 (chipmulties_11_cm_nx503), .A1 (
          chipmulties_11_cm_nx523)) ;
    aoi32 chipmulties_11_cm_ix524 (.Y (chipmulties_11_cm_nx523), .A0 (
          chipmulties_11_cm_nx52), .A1 (chipmulties_11_cm_nx54), .A2 (
          chipmulties_11_cm_nx28), .B0 (chipmulties_11_cm_nx46), .B1 (
          chipmulties_11_cm_nx68)) ;
    nor02 chipmulties_11_cm_ix53 (.Y (chipmulties_11_cm_nx52), .A0 (B_11__1), .A1 (
          chipmulties_11_cm_nx46)) ;
    nand02 chipmulties_11_cm_ix47 (.Y (chipmulties_11_cm_nx46), .A0 (A_11__0), .A1 (
           A_11__1)) ;
    nand02 chipmulties_11_cm_ix55 (.Y (chipmulties_11_cm_nx54), .A0 (
           chipmulties_11_cm_nx511), .A1 (chipmulties_11_cm_nx528)) ;
    inv01 chipmulties_11_cm_ix529 (.Y (chipmulties_11_cm_nx528), .A (B_11__4)) ;
    ao32 chipmulties_11_cm_ix69 (.Y (chipmulties_11_cm_nx68), .A0 (B_11__1), .A1 (
         A_11__0), .A2 (chipmulties_11_cm_nx62), .B0 (A_11__1), .B1 (
         chipmulties_11_cm_nx28)) ;
    aoi21 chipmulties_11_cm_ix63 (.Y (chipmulties_11_cm_nx62), .A0 (
          chipmulties_11_cm_nx511), .A1 (chipmulties_11_cm_nx528), .B0 (
          chipmulties_11_cm_nx508)) ;
    nor04 chipmulties_11_cm_ix109 (.Y (C_11__2), .A0 (chipmulties_11_cm_nx508), 
          .A1 (chipmulties_11_cm_nx533), .A2 (chipmulties_11_cm_nx535), .A3 (
          chipmulties_11_cm_nx537)) ;
    inv01 chipmulties_11_cm_ix534 (.Y (chipmulties_11_cm_nx533), .A (B_11__0)) ;
    nor03 chipmulties_11_cm_ix536 (.Y (chipmulties_11_cm_nx535), .A0 (A_11__0), 
          .A1 (A_11__1), .A2 (A_11__2)) ;
    ao22 chipmulties_11_cm_ix538 (.Y (chipmulties_11_cm_nx537), .A0 (
         chipmulties_11_cm_nx539), .A1 (chipmulties_11_cm_nx543), .B0 (
         chipmulties_11_cm_nx545), .B1 (chipmulties_11_cm_nx547)) ;
    oai21 chipmulties_11_cm_ix540 (.Y (chipmulties_11_cm_nx539), .A0 (A_11__2), 
          .A1 (B_11__1), .B0 (chipmulties_11_cm_nx541)) ;
    nor02 chipmulties_11_cm_ix542 (.Y (chipmulties_11_cm_nx541), .A0 (A_11__0), 
          .A1 (A_11__1)) ;
    xnor2 chipmulties_11_cm_ix544 (.Y (chipmulties_11_cm_nx543), .A0 (B_11__1), 
          .A1 (A_11__2)) ;
    oai22 chipmulties_11_cm_ix546 (.Y (chipmulties_11_cm_nx545), .A0 (
          chipmulties_11_cm_nx2), .A1 (chipmulties_11_cm_nx528), .B0 (
          chipmulties_11_cm_nx506), .B1 (A_11__4)) ;
    nand03 chipmulties_11_cm_ix548 (.Y (chipmulties_11_cm_nx547), .A0 (
           chipmulties_11_cm_nx2), .A1 (B_11__4), .A2 (chipmulties_11_cm_nx46)
           ) ;
    aoi21 chipmulties_11_cm_ix185 (.Y (C_11__3), .A0 (chipmulties_11_cm_nx550), 
          .A1 (chipmulties_11_cm_nx569), .B0 (chipmulties_11_cm_nx575)) ;
    oai21 chipmulties_11_cm_ix551 (.Y (chipmulties_11_cm_nx550), .A0 (
          chipmulties_11_cm_nx2), .A1 (A_11__1), .B0 (chipmulties_11_cm_nx178)
          ) ;
    oai22 chipmulties_11_cm_ix179 (.Y (chipmulties_11_cm_nx178), .A0 (
          chipmulties_11_cm_nx553), .A1 (chipmulties_11_cm_nx557), .B0 (
          chipmulties_11_cm_nx528), .B1 (chipmulties_11_cm_nx566)) ;
    aoi21 chipmulties_11_cm_ix554 (.Y (chipmulties_11_cm_nx553), .A0 (
          chipmulties_11_cm_nx555), .A1 (chipmulties_11_cm_nx46), .B0 (A_11__4)
          ) ;
    inv01 chipmulties_11_cm_ix556 (.Y (chipmulties_11_cm_nx555), .A (A_11__2)) ;
    nand02 chipmulties_11_cm_ix558 (.Y (chipmulties_11_cm_nx557), .A0 (
           chipmulties_11_cm_nx528), .A1 (chipmulties_11_cm_nx154)) ;
    oai21 chipmulties_11_cm_ix155 (.Y (chipmulties_11_cm_nx154), .A0 (
          chipmulties_11_cm_nx506), .A1 (A_11__0), .B0 (chipmulties_11_cm_nx560)
          ) ;
    aoi22 chipmulties_11_cm_ix561 (.Y (chipmulties_11_cm_nx560), .A0 (
          chipmulties_11_cm_nx562), .A1 (A_11__3), .B0 (chipmulties_11_cm_nx78)
          , .B1 (chipmulties_11_cm_nx130)) ;
    inv01 chipmulties_11_cm_ix563 (.Y (chipmulties_11_cm_nx562), .A (B_11__1)) ;
    aoi32 chipmulties_11_cm_ix567 (.Y (chipmulties_11_cm_nx566), .A0 (
          chipmulties_11_cm_nx164), .A1 (chipmulties_11_cm_nx78), .A2 (
          chipmulties_11_cm_nx130), .B0 (A_11__3), .B1 (chipmulties_11_cm_nx541)
          ) ;
    nand02 chipmulties_11_cm_ix165 (.Y (chipmulties_11_cm_nx164), .A0 (
           chipmulties_11_cm_nx555), .A1 (A_11__4)) ;
    or04 chipmulties_11_cm_ix570 (.Y (chipmulties_11_cm_nx569), .A0 (
         chipmulties_11_cm_nx528), .A1 (A_11__1), .A2 (chipmulties_11_cm_nx560)
         , .A3 (chipmulties_11_cm_nx571)) ;
    inv01 chipmulties_11_cm_ix574 (.Y (chipmulties_11_cm_nx573), .A (A_11__4)) ;
    nand03 chipmulties_11_cm_ix576 (.Y (chipmulties_11_cm_nx575), .A0 (
           chipmulties_11_cm_nx118), .A1 (B_11__0), .A2 (chipmulties_11_cm_nx18)
           ) ;
    nand03 chipmulties_11_cm_ix119 (.Y (chipmulties_11_cm_nx118), .A0 (B_11__4)
           , .A1 (A_11__2), .A2 (A_11__3)) ;
    nor02 chipmulties_11_cm_ix233 (.Y (C_11__4), .A0 (chipmulties_11_cm_nx575), 
          .A1 (chipmulties_11_cm_nx580)) ;
    aoi21 chipmulties_11_cm_ix581 (.Y (chipmulties_11_cm_nx580), .A0 (B_11__1), 
          .A1 (chipmulties_11_cm_nx192), .B0 (chipmulties_11_cm_nx228)) ;
    aoi21 chipmulties_11_cm_ix193 (.Y (chipmulties_11_cm_nx192), .A0 (
          chipmulties_11_cm_nx583), .A1 (B_11__4), .B0 (chipmulties_11_cm_nx22)
          ) ;
    oai33 chipmulties_11_cm_ix229 (.Y (chipmulties_11_cm_nx228), .A0 (
          chipmulties_11_cm_nx587), .A1 (chipmulties_11_cm_nx535), .A2 (
          chipmulties_11_cm_nx589), .B0 (B_11__1), .B1 (chipmulties_11_cm_nx573)
          , .B2 (chipmulties_11_cm_nx591)) ;
    aoi22 chipmulties_11_cm_ix588 (.Y (chipmulties_11_cm_nx587), .A0 (
          chipmulties_11_cm_nx562), .A1 (chipmulties_11_cm_nx571), .B0 (
          chipmulties_11_cm_nx573), .B1 (chipmulties_11_cm_nx130)) ;
    aoi21 chipmulties_11_cm_ix590 (.Y (chipmulties_11_cm_nx589), .A0 (A_11__2), 
          .A1 (A_11__1), .B0 (B_11__4)) ;
    oai21 chipmulties_11_cm_ix592 (.Y (chipmulties_11_cm_nx591), .A0 (
          chipmulties_11_cm_nx46), .A1 (chipmulties_11_cm_nx528), .B0 (A_11__3)
          ) ;
    inv01 chipmulties_11_cm_ix79 (.Y (chipmulties_11_cm_nx78), .A (
          chipmulties_11_cm_nx535)) ;
    inv01 chipmulties_11_cm_ix584 (.Y (chipmulties_11_cm_nx583), .A (
          chipmulties_11_cm_nx46)) ;
    inv01 chipmulties_11_cm_ix23 (.Y (chipmulties_11_cm_nx22), .A (
          chipmulties_11_cm_nx511)) ;
    inv01 chipmulties_11_cm_ix19 (.Y (chipmulties_11_cm_nx18), .A (
          chipmulties_11_cm_nx513)) ;
    inv01 chipmulties_11_cm_ix572 (.Y (chipmulties_11_cm_nx571), .A (
          chipmulties_11_cm_nx2)) ;
    nor02ii chipmulties_11_cm_ix512 (.Y (chipmulties_11_cm_nx511), .A0 (A_11__4)
            , .A1 (A_11__3)) ;
    and03 chipmulties_11_cm_ix519 (.Y (chipmulties_11_cm_nx518), .A0 (A_11__3), 
          .A1 (chipmulties_11_cm_nx573), .A2 (A_11__1)) ;
    nor02ii chipmulties_11_cm_ix131 (.Y (chipmulties_11_cm_nx130), .A0 (A_11__3)
            , .A1 (B_11__1)) ;
    nor04 chipmulties_10_cm_ix41 (.Y (C_10__0), .A0 (chipmulties_10_cm_nx501), .A1 (
          chipmulties_10_cm_nx503), .A2 (chipmulties_10_cm_nx508), .A3 (
          chipmulties_10_cm_nx518)) ;
    inv01 chipmulties_10_cm_ix502 (.Y (chipmulties_10_cm_nx501), .A (A_10__0)) ;
    oai21 chipmulties_10_cm_ix504 (.Y (chipmulties_10_cm_nx503), .A0 (
          chipmulties_10_cm_nx2), .A1 (A_10__2), .B0 (B_10__0)) ;
    nand02 chipmulties_10_cm_ix3 (.Y (chipmulties_10_cm_nx2), .A0 (
           chipmulties_10_cm_nx506), .A1 (A_10__4)) ;
    inv01 chipmulties_10_cm_ix507 (.Y (chipmulties_10_cm_nx506), .A (A_10__3)) ;
    oai21 chipmulties_10_cm_ix509 (.Y (chipmulties_10_cm_nx508), .A0 (
          chipmulties_10_cm_nx2), .A1 (A_10__1), .B0 (chipmulties_10_cm_nx28)) ;
    aoi21 chipmulties_10_cm_ix29 (.Y (chipmulties_10_cm_nx28), .A0 (
          chipmulties_10_cm_nx511), .A1 (A_10__2), .B0 (chipmulties_10_cm_nx513)
          ) ;
    nand03 chipmulties_10_cm_ix514 (.Y (chipmulties_10_cm_nx513), .A0 (
           chipmulties_10_cm_nx10), .A1 (chipmulties_10_cm_nx12), .A2 (
           chipmulties_10_cm_nx14)) ;
    xnor2 chipmulties_10_cm_ix11 (.Y (chipmulties_10_cm_nx10), .A0 (B_10__3), .A1 (
          B_10__4)) ;
    xnor2 chipmulties_10_cm_ix13 (.Y (chipmulties_10_cm_nx12), .A0 (B_10__2), .A1 (
          B_10__1)) ;
    xnor2 chipmulties_10_cm_ix15 (.Y (chipmulties_10_cm_nx14), .A0 (B_10__3), .A1 (
          B_10__2)) ;
    nor02 chipmulties_10_cm_ix75 (.Y (C_10__1), .A0 (chipmulties_10_cm_nx503), .A1 (
          chipmulties_10_cm_nx523)) ;
    aoi32 chipmulties_10_cm_ix524 (.Y (chipmulties_10_cm_nx523), .A0 (
          chipmulties_10_cm_nx52), .A1 (chipmulties_10_cm_nx54), .A2 (
          chipmulties_10_cm_nx28), .B0 (chipmulties_10_cm_nx46), .B1 (
          chipmulties_10_cm_nx68)) ;
    nor02 chipmulties_10_cm_ix53 (.Y (chipmulties_10_cm_nx52), .A0 (B_10__1), .A1 (
          chipmulties_10_cm_nx46)) ;
    nand02 chipmulties_10_cm_ix47 (.Y (chipmulties_10_cm_nx46), .A0 (A_10__0), .A1 (
           A_10__1)) ;
    nand02 chipmulties_10_cm_ix55 (.Y (chipmulties_10_cm_nx54), .A0 (
           chipmulties_10_cm_nx511), .A1 (chipmulties_10_cm_nx528)) ;
    inv01 chipmulties_10_cm_ix529 (.Y (chipmulties_10_cm_nx528), .A (B_10__4)) ;
    ao32 chipmulties_10_cm_ix69 (.Y (chipmulties_10_cm_nx68), .A0 (B_10__1), .A1 (
         A_10__0), .A2 (chipmulties_10_cm_nx62), .B0 (A_10__1), .B1 (
         chipmulties_10_cm_nx28)) ;
    aoi21 chipmulties_10_cm_ix63 (.Y (chipmulties_10_cm_nx62), .A0 (
          chipmulties_10_cm_nx511), .A1 (chipmulties_10_cm_nx528), .B0 (
          chipmulties_10_cm_nx508)) ;
    nor04 chipmulties_10_cm_ix109 (.Y (C_10__2), .A0 (chipmulties_10_cm_nx508), 
          .A1 (chipmulties_10_cm_nx533), .A2 (chipmulties_10_cm_nx535), .A3 (
          chipmulties_10_cm_nx537)) ;
    inv01 chipmulties_10_cm_ix534 (.Y (chipmulties_10_cm_nx533), .A (B_10__0)) ;
    nor03 chipmulties_10_cm_ix536 (.Y (chipmulties_10_cm_nx535), .A0 (A_10__0), 
          .A1 (A_10__1), .A2 (A_10__2)) ;
    ao22 chipmulties_10_cm_ix538 (.Y (chipmulties_10_cm_nx537), .A0 (
         chipmulties_10_cm_nx539), .A1 (chipmulties_10_cm_nx543), .B0 (
         chipmulties_10_cm_nx545), .B1 (chipmulties_10_cm_nx547)) ;
    oai21 chipmulties_10_cm_ix540 (.Y (chipmulties_10_cm_nx539), .A0 (A_10__2), 
          .A1 (B_10__1), .B0 (chipmulties_10_cm_nx541)) ;
    nor02 chipmulties_10_cm_ix542 (.Y (chipmulties_10_cm_nx541), .A0 (A_10__0), 
          .A1 (A_10__1)) ;
    xnor2 chipmulties_10_cm_ix544 (.Y (chipmulties_10_cm_nx543), .A0 (B_10__1), 
          .A1 (A_10__2)) ;
    oai22 chipmulties_10_cm_ix546 (.Y (chipmulties_10_cm_nx545), .A0 (
          chipmulties_10_cm_nx2), .A1 (chipmulties_10_cm_nx528), .B0 (
          chipmulties_10_cm_nx506), .B1 (A_10__4)) ;
    nand03 chipmulties_10_cm_ix548 (.Y (chipmulties_10_cm_nx547), .A0 (
           chipmulties_10_cm_nx2), .A1 (B_10__4), .A2 (chipmulties_10_cm_nx46)
           ) ;
    aoi21 chipmulties_10_cm_ix185 (.Y (C_10__3), .A0 (chipmulties_10_cm_nx550), 
          .A1 (chipmulties_10_cm_nx569), .B0 (chipmulties_10_cm_nx575)) ;
    oai21 chipmulties_10_cm_ix551 (.Y (chipmulties_10_cm_nx550), .A0 (
          chipmulties_10_cm_nx2), .A1 (A_10__1), .B0 (chipmulties_10_cm_nx178)
          ) ;
    oai22 chipmulties_10_cm_ix179 (.Y (chipmulties_10_cm_nx178), .A0 (
          chipmulties_10_cm_nx553), .A1 (chipmulties_10_cm_nx557), .B0 (
          chipmulties_10_cm_nx528), .B1 (chipmulties_10_cm_nx566)) ;
    aoi21 chipmulties_10_cm_ix554 (.Y (chipmulties_10_cm_nx553), .A0 (
          chipmulties_10_cm_nx555), .A1 (chipmulties_10_cm_nx46), .B0 (A_10__4)
          ) ;
    inv01 chipmulties_10_cm_ix556 (.Y (chipmulties_10_cm_nx555), .A (A_10__2)) ;
    nand02 chipmulties_10_cm_ix558 (.Y (chipmulties_10_cm_nx557), .A0 (
           chipmulties_10_cm_nx528), .A1 (chipmulties_10_cm_nx154)) ;
    oai21 chipmulties_10_cm_ix155 (.Y (chipmulties_10_cm_nx154), .A0 (
          chipmulties_10_cm_nx506), .A1 (A_10__0), .B0 (chipmulties_10_cm_nx560)
          ) ;
    aoi22 chipmulties_10_cm_ix561 (.Y (chipmulties_10_cm_nx560), .A0 (
          chipmulties_10_cm_nx562), .A1 (A_10__3), .B0 (chipmulties_10_cm_nx78)
          , .B1 (chipmulties_10_cm_nx130)) ;
    inv01 chipmulties_10_cm_ix563 (.Y (chipmulties_10_cm_nx562), .A (B_10__1)) ;
    aoi32 chipmulties_10_cm_ix567 (.Y (chipmulties_10_cm_nx566), .A0 (
          chipmulties_10_cm_nx164), .A1 (chipmulties_10_cm_nx78), .A2 (
          chipmulties_10_cm_nx130), .B0 (A_10__3), .B1 (chipmulties_10_cm_nx541)
          ) ;
    nand02 chipmulties_10_cm_ix165 (.Y (chipmulties_10_cm_nx164), .A0 (
           chipmulties_10_cm_nx555), .A1 (A_10__4)) ;
    or04 chipmulties_10_cm_ix570 (.Y (chipmulties_10_cm_nx569), .A0 (
         chipmulties_10_cm_nx528), .A1 (A_10__1), .A2 (chipmulties_10_cm_nx560)
         , .A3 (chipmulties_10_cm_nx571)) ;
    inv01 chipmulties_10_cm_ix574 (.Y (chipmulties_10_cm_nx573), .A (A_10__4)) ;
    nand03 chipmulties_10_cm_ix576 (.Y (chipmulties_10_cm_nx575), .A0 (
           chipmulties_10_cm_nx118), .A1 (B_10__0), .A2 (chipmulties_10_cm_nx18)
           ) ;
    nand03 chipmulties_10_cm_ix119 (.Y (chipmulties_10_cm_nx118), .A0 (B_10__4)
           , .A1 (A_10__2), .A2 (A_10__3)) ;
    nor02 chipmulties_10_cm_ix233 (.Y (C_10__4), .A0 (chipmulties_10_cm_nx575), 
          .A1 (chipmulties_10_cm_nx580)) ;
    aoi21 chipmulties_10_cm_ix581 (.Y (chipmulties_10_cm_nx580), .A0 (B_10__1), 
          .A1 (chipmulties_10_cm_nx192), .B0 (chipmulties_10_cm_nx228)) ;
    aoi21 chipmulties_10_cm_ix193 (.Y (chipmulties_10_cm_nx192), .A0 (
          chipmulties_10_cm_nx583), .A1 (B_10__4), .B0 (chipmulties_10_cm_nx22)
          ) ;
    oai33 chipmulties_10_cm_ix229 (.Y (chipmulties_10_cm_nx228), .A0 (
          chipmulties_10_cm_nx587), .A1 (chipmulties_10_cm_nx535), .A2 (
          chipmulties_10_cm_nx589), .B0 (B_10__1), .B1 (chipmulties_10_cm_nx573)
          , .B2 (chipmulties_10_cm_nx591)) ;
    aoi22 chipmulties_10_cm_ix588 (.Y (chipmulties_10_cm_nx587), .A0 (
          chipmulties_10_cm_nx562), .A1 (chipmulties_10_cm_nx571), .B0 (
          chipmulties_10_cm_nx573), .B1 (chipmulties_10_cm_nx130)) ;
    aoi21 chipmulties_10_cm_ix590 (.Y (chipmulties_10_cm_nx589), .A0 (A_10__2), 
          .A1 (A_10__1), .B0 (B_10__4)) ;
    oai21 chipmulties_10_cm_ix592 (.Y (chipmulties_10_cm_nx591), .A0 (
          chipmulties_10_cm_nx46), .A1 (chipmulties_10_cm_nx528), .B0 (A_10__3)
          ) ;
    inv01 chipmulties_10_cm_ix79 (.Y (chipmulties_10_cm_nx78), .A (
          chipmulties_10_cm_nx535)) ;
    inv01 chipmulties_10_cm_ix584 (.Y (chipmulties_10_cm_nx583), .A (
          chipmulties_10_cm_nx46)) ;
    inv01 chipmulties_10_cm_ix23 (.Y (chipmulties_10_cm_nx22), .A (
          chipmulties_10_cm_nx511)) ;
    inv01 chipmulties_10_cm_ix19 (.Y (chipmulties_10_cm_nx18), .A (
          chipmulties_10_cm_nx513)) ;
    inv01 chipmulties_10_cm_ix572 (.Y (chipmulties_10_cm_nx571), .A (
          chipmulties_10_cm_nx2)) ;
    nor02ii chipmulties_10_cm_ix512 (.Y (chipmulties_10_cm_nx511), .A0 (A_10__4)
            , .A1 (A_10__3)) ;
    and03 chipmulties_10_cm_ix519 (.Y (chipmulties_10_cm_nx518), .A0 (A_10__3), 
          .A1 (chipmulties_10_cm_nx573), .A2 (A_10__1)) ;
    nor02ii chipmulties_10_cm_ix131 (.Y (chipmulties_10_cm_nx130), .A0 (A_10__3)
            , .A1 (B_10__1)) ;
    nor04 chipmulties_9_cm_ix41 (.Y (C_9__0), .A0 (chipmulties_9_cm_nx501), .A1 (
          chipmulties_9_cm_nx503), .A2 (chipmulties_9_cm_nx508), .A3 (
          chipmulties_9_cm_nx518)) ;
    inv01 chipmulties_9_cm_ix502 (.Y (chipmulties_9_cm_nx501), .A (A_9__0)) ;
    oai21 chipmulties_9_cm_ix504 (.Y (chipmulties_9_cm_nx503), .A0 (
          chipmulties_9_cm_nx2), .A1 (A_9__2), .B0 (B_9__0)) ;
    nand02 chipmulties_9_cm_ix3 (.Y (chipmulties_9_cm_nx2), .A0 (
           chipmulties_9_cm_nx506), .A1 (A_9__4)) ;
    inv01 chipmulties_9_cm_ix507 (.Y (chipmulties_9_cm_nx506), .A (A_9__3)) ;
    oai21 chipmulties_9_cm_ix509 (.Y (chipmulties_9_cm_nx508), .A0 (
          chipmulties_9_cm_nx2), .A1 (A_9__1), .B0 (chipmulties_9_cm_nx28)) ;
    aoi21 chipmulties_9_cm_ix29 (.Y (chipmulties_9_cm_nx28), .A0 (
          chipmulties_9_cm_nx511), .A1 (A_9__2), .B0 (chipmulties_9_cm_nx513)) ;
    nand03 chipmulties_9_cm_ix514 (.Y (chipmulties_9_cm_nx513), .A0 (
           chipmulties_9_cm_nx10), .A1 (chipmulties_9_cm_nx12), .A2 (
           chipmulties_9_cm_nx14)) ;
    xnor2 chipmulties_9_cm_ix11 (.Y (chipmulties_9_cm_nx10), .A0 (B_9__3), .A1 (
          B_9__4)) ;
    xnor2 chipmulties_9_cm_ix13 (.Y (chipmulties_9_cm_nx12), .A0 (B_9__2), .A1 (
          B_9__1)) ;
    xnor2 chipmulties_9_cm_ix15 (.Y (chipmulties_9_cm_nx14), .A0 (B_9__3), .A1 (
          B_9__2)) ;
    nor02 chipmulties_9_cm_ix75 (.Y (C_9__1), .A0 (chipmulties_9_cm_nx503), .A1 (
          chipmulties_9_cm_nx523)) ;
    aoi32 chipmulties_9_cm_ix524 (.Y (chipmulties_9_cm_nx523), .A0 (
          chipmulties_9_cm_nx52), .A1 (chipmulties_9_cm_nx54), .A2 (
          chipmulties_9_cm_nx28), .B0 (chipmulties_9_cm_nx46), .B1 (
          chipmulties_9_cm_nx68)) ;
    nor02 chipmulties_9_cm_ix53 (.Y (chipmulties_9_cm_nx52), .A0 (B_9__1), .A1 (
          chipmulties_9_cm_nx46)) ;
    nand02 chipmulties_9_cm_ix47 (.Y (chipmulties_9_cm_nx46), .A0 (A_9__0), .A1 (
           A_9__1)) ;
    nand02 chipmulties_9_cm_ix55 (.Y (chipmulties_9_cm_nx54), .A0 (
           chipmulties_9_cm_nx511), .A1 (chipmulties_9_cm_nx528)) ;
    inv01 chipmulties_9_cm_ix529 (.Y (chipmulties_9_cm_nx528), .A (B_9__4)) ;
    ao32 chipmulties_9_cm_ix69 (.Y (chipmulties_9_cm_nx68), .A0 (B_9__1), .A1 (
         A_9__0), .A2 (chipmulties_9_cm_nx62), .B0 (A_9__1), .B1 (
         chipmulties_9_cm_nx28)) ;
    aoi21 chipmulties_9_cm_ix63 (.Y (chipmulties_9_cm_nx62), .A0 (
          chipmulties_9_cm_nx511), .A1 (chipmulties_9_cm_nx528), .B0 (
          chipmulties_9_cm_nx508)) ;
    nor04 chipmulties_9_cm_ix109 (.Y (C_9__2), .A0 (chipmulties_9_cm_nx508), .A1 (
          chipmulties_9_cm_nx533), .A2 (chipmulties_9_cm_nx535), .A3 (
          chipmulties_9_cm_nx537)) ;
    inv01 chipmulties_9_cm_ix534 (.Y (chipmulties_9_cm_nx533), .A (B_9__0)) ;
    nor03 chipmulties_9_cm_ix536 (.Y (chipmulties_9_cm_nx535), .A0 (A_9__0), .A1 (
          A_9__1), .A2 (A_9__2)) ;
    ao22 chipmulties_9_cm_ix538 (.Y (chipmulties_9_cm_nx537), .A0 (
         chipmulties_9_cm_nx539), .A1 (chipmulties_9_cm_nx543), .B0 (
         chipmulties_9_cm_nx545), .B1 (chipmulties_9_cm_nx547)) ;
    oai21 chipmulties_9_cm_ix540 (.Y (chipmulties_9_cm_nx539), .A0 (A_9__2), .A1 (
          B_9__1), .B0 (chipmulties_9_cm_nx541)) ;
    nor02 chipmulties_9_cm_ix542 (.Y (chipmulties_9_cm_nx541), .A0 (A_9__0), .A1 (
          A_9__1)) ;
    xnor2 chipmulties_9_cm_ix544 (.Y (chipmulties_9_cm_nx543), .A0 (B_9__1), .A1 (
          A_9__2)) ;
    oai22 chipmulties_9_cm_ix546 (.Y (chipmulties_9_cm_nx545), .A0 (
          chipmulties_9_cm_nx2), .A1 (chipmulties_9_cm_nx528), .B0 (
          chipmulties_9_cm_nx506), .B1 (A_9__4)) ;
    nand03 chipmulties_9_cm_ix548 (.Y (chipmulties_9_cm_nx547), .A0 (
           chipmulties_9_cm_nx2), .A1 (B_9__4), .A2 (chipmulties_9_cm_nx46)) ;
    aoi21 chipmulties_9_cm_ix185 (.Y (C_9__3), .A0 (chipmulties_9_cm_nx550), .A1 (
          chipmulties_9_cm_nx569), .B0 (chipmulties_9_cm_nx575)) ;
    oai21 chipmulties_9_cm_ix551 (.Y (chipmulties_9_cm_nx550), .A0 (
          chipmulties_9_cm_nx2), .A1 (A_9__1), .B0 (chipmulties_9_cm_nx178)) ;
    oai22 chipmulties_9_cm_ix179 (.Y (chipmulties_9_cm_nx178), .A0 (
          chipmulties_9_cm_nx553), .A1 (chipmulties_9_cm_nx557), .B0 (
          chipmulties_9_cm_nx528), .B1 (chipmulties_9_cm_nx566)) ;
    aoi21 chipmulties_9_cm_ix554 (.Y (chipmulties_9_cm_nx553), .A0 (
          chipmulties_9_cm_nx555), .A1 (chipmulties_9_cm_nx46), .B0 (A_9__4)) ;
    inv01 chipmulties_9_cm_ix556 (.Y (chipmulties_9_cm_nx555), .A (A_9__2)) ;
    nand02 chipmulties_9_cm_ix558 (.Y (chipmulties_9_cm_nx557), .A0 (
           chipmulties_9_cm_nx528), .A1 (chipmulties_9_cm_nx154)) ;
    oai21 chipmulties_9_cm_ix155 (.Y (chipmulties_9_cm_nx154), .A0 (
          chipmulties_9_cm_nx506), .A1 (A_9__0), .B0 (chipmulties_9_cm_nx560)) ;
    aoi22 chipmulties_9_cm_ix561 (.Y (chipmulties_9_cm_nx560), .A0 (
          chipmulties_9_cm_nx562), .A1 (A_9__3), .B0 (chipmulties_9_cm_nx78), .B1 (
          chipmulties_9_cm_nx130)) ;
    inv01 chipmulties_9_cm_ix563 (.Y (chipmulties_9_cm_nx562), .A (B_9__1)) ;
    aoi32 chipmulties_9_cm_ix567 (.Y (chipmulties_9_cm_nx566), .A0 (
          chipmulties_9_cm_nx164), .A1 (chipmulties_9_cm_nx78), .A2 (
          chipmulties_9_cm_nx130), .B0 (A_9__3), .B1 (chipmulties_9_cm_nx541)) ;
    nand02 chipmulties_9_cm_ix165 (.Y (chipmulties_9_cm_nx164), .A0 (
           chipmulties_9_cm_nx555), .A1 (A_9__4)) ;
    or04 chipmulties_9_cm_ix570 (.Y (chipmulties_9_cm_nx569), .A0 (
         chipmulties_9_cm_nx528), .A1 (A_9__1), .A2 (chipmulties_9_cm_nx560), .A3 (
         chipmulties_9_cm_nx571)) ;
    inv01 chipmulties_9_cm_ix574 (.Y (chipmulties_9_cm_nx573), .A (A_9__4)) ;
    nand03 chipmulties_9_cm_ix576 (.Y (chipmulties_9_cm_nx575), .A0 (
           chipmulties_9_cm_nx118), .A1 (B_9__0), .A2 (chipmulties_9_cm_nx18)) ;
    nand03 chipmulties_9_cm_ix119 (.Y (chipmulties_9_cm_nx118), .A0 (B_9__4), .A1 (
           A_9__2), .A2 (A_9__3)) ;
    nor02 chipmulties_9_cm_ix233 (.Y (C_9__4), .A0 (chipmulties_9_cm_nx575), .A1 (
          chipmulties_9_cm_nx580)) ;
    aoi21 chipmulties_9_cm_ix581 (.Y (chipmulties_9_cm_nx580), .A0 (B_9__1), .A1 (
          chipmulties_9_cm_nx192), .B0 (chipmulties_9_cm_nx228)) ;
    aoi21 chipmulties_9_cm_ix193 (.Y (chipmulties_9_cm_nx192), .A0 (
          chipmulties_9_cm_nx583), .A1 (B_9__4), .B0 (chipmulties_9_cm_nx22)) ;
    oai33 chipmulties_9_cm_ix229 (.Y (chipmulties_9_cm_nx228), .A0 (
          chipmulties_9_cm_nx587), .A1 (chipmulties_9_cm_nx535), .A2 (
          chipmulties_9_cm_nx589), .B0 (B_9__1), .B1 (chipmulties_9_cm_nx573), .B2 (
          chipmulties_9_cm_nx591)) ;
    aoi22 chipmulties_9_cm_ix588 (.Y (chipmulties_9_cm_nx587), .A0 (
          chipmulties_9_cm_nx562), .A1 (chipmulties_9_cm_nx571), .B0 (
          chipmulties_9_cm_nx573), .B1 (chipmulties_9_cm_nx130)) ;
    aoi21 chipmulties_9_cm_ix590 (.Y (chipmulties_9_cm_nx589), .A0 (A_9__2), .A1 (
          A_9__1), .B0 (B_9__4)) ;
    oai21 chipmulties_9_cm_ix592 (.Y (chipmulties_9_cm_nx591), .A0 (
          chipmulties_9_cm_nx46), .A1 (chipmulties_9_cm_nx528), .B0 (A_9__3)) ;
    inv01 chipmulties_9_cm_ix79 (.Y (chipmulties_9_cm_nx78), .A (
          chipmulties_9_cm_nx535)) ;
    inv01 chipmulties_9_cm_ix584 (.Y (chipmulties_9_cm_nx583), .A (
          chipmulties_9_cm_nx46)) ;
    inv01 chipmulties_9_cm_ix23 (.Y (chipmulties_9_cm_nx22), .A (
          chipmulties_9_cm_nx511)) ;
    inv01 chipmulties_9_cm_ix19 (.Y (chipmulties_9_cm_nx18), .A (
          chipmulties_9_cm_nx513)) ;
    inv01 chipmulties_9_cm_ix572 (.Y (chipmulties_9_cm_nx571), .A (
          chipmulties_9_cm_nx2)) ;
    nor02ii chipmulties_9_cm_ix512 (.Y (chipmulties_9_cm_nx511), .A0 (A_9__4), .A1 (
            A_9__3)) ;
    and03 chipmulties_9_cm_ix519 (.Y (chipmulties_9_cm_nx518), .A0 (A_9__3), .A1 (
          chipmulties_9_cm_nx573), .A2 (A_9__1)) ;
    nor02ii chipmulties_9_cm_ix131 (.Y (chipmulties_9_cm_nx130), .A0 (A_9__3), .A1 (
            B_9__1)) ;
    nor04 chipmulties_8_cm_ix41 (.Y (C_8__0), .A0 (chipmulties_8_cm_nx501), .A1 (
          chipmulties_8_cm_nx503), .A2 (chipmulties_8_cm_nx508), .A3 (
          chipmulties_8_cm_nx518)) ;
    inv01 chipmulties_8_cm_ix502 (.Y (chipmulties_8_cm_nx501), .A (A_8__0)) ;
    oai21 chipmulties_8_cm_ix504 (.Y (chipmulties_8_cm_nx503), .A0 (
          chipmulties_8_cm_nx2), .A1 (A_8__2), .B0 (B_8__0)) ;
    nand02 chipmulties_8_cm_ix3 (.Y (chipmulties_8_cm_nx2), .A0 (
           chipmulties_8_cm_nx506), .A1 (A_8__4)) ;
    inv01 chipmulties_8_cm_ix507 (.Y (chipmulties_8_cm_nx506), .A (A_8__3)) ;
    oai21 chipmulties_8_cm_ix509 (.Y (chipmulties_8_cm_nx508), .A0 (
          chipmulties_8_cm_nx2), .A1 (A_8__1), .B0 (chipmulties_8_cm_nx28)) ;
    aoi21 chipmulties_8_cm_ix29 (.Y (chipmulties_8_cm_nx28), .A0 (
          chipmulties_8_cm_nx511), .A1 (A_8__2), .B0 (chipmulties_8_cm_nx513)) ;
    nand03 chipmulties_8_cm_ix514 (.Y (chipmulties_8_cm_nx513), .A0 (
           chipmulties_8_cm_nx10), .A1 (chipmulties_8_cm_nx12), .A2 (
           chipmulties_8_cm_nx14)) ;
    xnor2 chipmulties_8_cm_ix11 (.Y (chipmulties_8_cm_nx10), .A0 (B_8__3), .A1 (
          B_8__4)) ;
    xnor2 chipmulties_8_cm_ix13 (.Y (chipmulties_8_cm_nx12), .A0 (B_8__2), .A1 (
          B_8__1)) ;
    xnor2 chipmulties_8_cm_ix15 (.Y (chipmulties_8_cm_nx14), .A0 (B_8__3), .A1 (
          B_8__2)) ;
    nor02 chipmulties_8_cm_ix75 (.Y (C_8__1), .A0 (chipmulties_8_cm_nx503), .A1 (
          chipmulties_8_cm_nx523)) ;
    aoi32 chipmulties_8_cm_ix524 (.Y (chipmulties_8_cm_nx523), .A0 (
          chipmulties_8_cm_nx52), .A1 (chipmulties_8_cm_nx54), .A2 (
          chipmulties_8_cm_nx28), .B0 (chipmulties_8_cm_nx46), .B1 (
          chipmulties_8_cm_nx68)) ;
    nor02 chipmulties_8_cm_ix53 (.Y (chipmulties_8_cm_nx52), .A0 (B_8__1), .A1 (
          chipmulties_8_cm_nx46)) ;
    nand02 chipmulties_8_cm_ix47 (.Y (chipmulties_8_cm_nx46), .A0 (A_8__0), .A1 (
           A_8__1)) ;
    nand02 chipmulties_8_cm_ix55 (.Y (chipmulties_8_cm_nx54), .A0 (
           chipmulties_8_cm_nx511), .A1 (chipmulties_8_cm_nx528)) ;
    inv01 chipmulties_8_cm_ix529 (.Y (chipmulties_8_cm_nx528), .A (B_8__4)) ;
    ao32 chipmulties_8_cm_ix69 (.Y (chipmulties_8_cm_nx68), .A0 (B_8__1), .A1 (
         A_8__0), .A2 (chipmulties_8_cm_nx62), .B0 (A_8__1), .B1 (
         chipmulties_8_cm_nx28)) ;
    aoi21 chipmulties_8_cm_ix63 (.Y (chipmulties_8_cm_nx62), .A0 (
          chipmulties_8_cm_nx511), .A1 (chipmulties_8_cm_nx528), .B0 (
          chipmulties_8_cm_nx508)) ;
    nor04 chipmulties_8_cm_ix109 (.Y (C_8__2), .A0 (chipmulties_8_cm_nx508), .A1 (
          chipmulties_8_cm_nx533), .A2 (chipmulties_8_cm_nx535), .A3 (
          chipmulties_8_cm_nx537)) ;
    inv01 chipmulties_8_cm_ix534 (.Y (chipmulties_8_cm_nx533), .A (B_8__0)) ;
    nor03 chipmulties_8_cm_ix536 (.Y (chipmulties_8_cm_nx535), .A0 (A_8__0), .A1 (
          A_8__1), .A2 (A_8__2)) ;
    ao22 chipmulties_8_cm_ix538 (.Y (chipmulties_8_cm_nx537), .A0 (
         chipmulties_8_cm_nx539), .A1 (chipmulties_8_cm_nx543), .B0 (
         chipmulties_8_cm_nx545), .B1 (chipmulties_8_cm_nx547)) ;
    oai21 chipmulties_8_cm_ix540 (.Y (chipmulties_8_cm_nx539), .A0 (A_8__2), .A1 (
          B_8__1), .B0 (chipmulties_8_cm_nx541)) ;
    nor02 chipmulties_8_cm_ix542 (.Y (chipmulties_8_cm_nx541), .A0 (A_8__0), .A1 (
          A_8__1)) ;
    xnor2 chipmulties_8_cm_ix544 (.Y (chipmulties_8_cm_nx543), .A0 (B_8__1), .A1 (
          A_8__2)) ;
    oai22 chipmulties_8_cm_ix546 (.Y (chipmulties_8_cm_nx545), .A0 (
          chipmulties_8_cm_nx2), .A1 (chipmulties_8_cm_nx528), .B0 (
          chipmulties_8_cm_nx506), .B1 (A_8__4)) ;
    nand03 chipmulties_8_cm_ix548 (.Y (chipmulties_8_cm_nx547), .A0 (
           chipmulties_8_cm_nx2), .A1 (B_8__4), .A2 (chipmulties_8_cm_nx46)) ;
    aoi21 chipmulties_8_cm_ix185 (.Y (C_8__3), .A0 (chipmulties_8_cm_nx550), .A1 (
          chipmulties_8_cm_nx569), .B0 (chipmulties_8_cm_nx575)) ;
    oai21 chipmulties_8_cm_ix551 (.Y (chipmulties_8_cm_nx550), .A0 (
          chipmulties_8_cm_nx2), .A1 (A_8__1), .B0 (chipmulties_8_cm_nx178)) ;
    oai22 chipmulties_8_cm_ix179 (.Y (chipmulties_8_cm_nx178), .A0 (
          chipmulties_8_cm_nx553), .A1 (chipmulties_8_cm_nx557), .B0 (
          chipmulties_8_cm_nx528), .B1 (chipmulties_8_cm_nx566)) ;
    aoi21 chipmulties_8_cm_ix554 (.Y (chipmulties_8_cm_nx553), .A0 (
          chipmulties_8_cm_nx555), .A1 (chipmulties_8_cm_nx46), .B0 (A_8__4)) ;
    inv01 chipmulties_8_cm_ix556 (.Y (chipmulties_8_cm_nx555), .A (A_8__2)) ;
    nand02 chipmulties_8_cm_ix558 (.Y (chipmulties_8_cm_nx557), .A0 (
           chipmulties_8_cm_nx528), .A1 (chipmulties_8_cm_nx154)) ;
    oai21 chipmulties_8_cm_ix155 (.Y (chipmulties_8_cm_nx154), .A0 (
          chipmulties_8_cm_nx506), .A1 (A_8__0), .B0 (chipmulties_8_cm_nx560)) ;
    aoi22 chipmulties_8_cm_ix561 (.Y (chipmulties_8_cm_nx560), .A0 (
          chipmulties_8_cm_nx562), .A1 (A_8__3), .B0 (chipmulties_8_cm_nx78), .B1 (
          chipmulties_8_cm_nx130)) ;
    inv01 chipmulties_8_cm_ix563 (.Y (chipmulties_8_cm_nx562), .A (B_8__1)) ;
    aoi32 chipmulties_8_cm_ix567 (.Y (chipmulties_8_cm_nx566), .A0 (
          chipmulties_8_cm_nx164), .A1 (chipmulties_8_cm_nx78), .A2 (
          chipmulties_8_cm_nx130), .B0 (A_8__3), .B1 (chipmulties_8_cm_nx541)) ;
    nand02 chipmulties_8_cm_ix165 (.Y (chipmulties_8_cm_nx164), .A0 (
           chipmulties_8_cm_nx555), .A1 (A_8__4)) ;
    or04 chipmulties_8_cm_ix570 (.Y (chipmulties_8_cm_nx569), .A0 (
         chipmulties_8_cm_nx528), .A1 (A_8__1), .A2 (chipmulties_8_cm_nx560), .A3 (
         chipmulties_8_cm_nx571)) ;
    inv01 chipmulties_8_cm_ix574 (.Y (chipmulties_8_cm_nx573), .A (A_8__4)) ;
    nand03 chipmulties_8_cm_ix576 (.Y (chipmulties_8_cm_nx575), .A0 (
           chipmulties_8_cm_nx118), .A1 (B_8__0), .A2 (chipmulties_8_cm_nx18)) ;
    nand03 chipmulties_8_cm_ix119 (.Y (chipmulties_8_cm_nx118), .A0 (B_8__4), .A1 (
           A_8__2), .A2 (A_8__3)) ;
    nor02 chipmulties_8_cm_ix233 (.Y (C_8__4), .A0 (chipmulties_8_cm_nx575), .A1 (
          chipmulties_8_cm_nx580)) ;
    aoi21 chipmulties_8_cm_ix581 (.Y (chipmulties_8_cm_nx580), .A0 (B_8__1), .A1 (
          chipmulties_8_cm_nx192), .B0 (chipmulties_8_cm_nx228)) ;
    aoi21 chipmulties_8_cm_ix193 (.Y (chipmulties_8_cm_nx192), .A0 (
          chipmulties_8_cm_nx583), .A1 (B_8__4), .B0 (chipmulties_8_cm_nx22)) ;
    oai33 chipmulties_8_cm_ix229 (.Y (chipmulties_8_cm_nx228), .A0 (
          chipmulties_8_cm_nx587), .A1 (chipmulties_8_cm_nx535), .A2 (
          chipmulties_8_cm_nx589), .B0 (B_8__1), .B1 (chipmulties_8_cm_nx573), .B2 (
          chipmulties_8_cm_nx591)) ;
    aoi22 chipmulties_8_cm_ix588 (.Y (chipmulties_8_cm_nx587), .A0 (
          chipmulties_8_cm_nx562), .A1 (chipmulties_8_cm_nx571), .B0 (
          chipmulties_8_cm_nx573), .B1 (chipmulties_8_cm_nx130)) ;
    aoi21 chipmulties_8_cm_ix590 (.Y (chipmulties_8_cm_nx589), .A0 (A_8__2), .A1 (
          A_8__1), .B0 (B_8__4)) ;
    oai21 chipmulties_8_cm_ix592 (.Y (chipmulties_8_cm_nx591), .A0 (
          chipmulties_8_cm_nx46), .A1 (chipmulties_8_cm_nx528), .B0 (A_8__3)) ;
    inv01 chipmulties_8_cm_ix79 (.Y (chipmulties_8_cm_nx78), .A (
          chipmulties_8_cm_nx535)) ;
    inv01 chipmulties_8_cm_ix584 (.Y (chipmulties_8_cm_nx583), .A (
          chipmulties_8_cm_nx46)) ;
    inv01 chipmulties_8_cm_ix23 (.Y (chipmulties_8_cm_nx22), .A (
          chipmulties_8_cm_nx511)) ;
    inv01 chipmulties_8_cm_ix19 (.Y (chipmulties_8_cm_nx18), .A (
          chipmulties_8_cm_nx513)) ;
    inv01 chipmulties_8_cm_ix572 (.Y (chipmulties_8_cm_nx571), .A (
          chipmulties_8_cm_nx2)) ;
    nor02ii chipmulties_8_cm_ix512 (.Y (chipmulties_8_cm_nx511), .A0 (A_8__4), .A1 (
            A_8__3)) ;
    and03 chipmulties_8_cm_ix519 (.Y (chipmulties_8_cm_nx518), .A0 (A_8__3), .A1 (
          chipmulties_8_cm_nx573), .A2 (A_8__1)) ;
    nor02ii chipmulties_8_cm_ix131 (.Y (chipmulties_8_cm_nx130), .A0 (A_8__3), .A1 (
            B_8__1)) ;
    nor04 chipmulties_7_cm_ix41 (.Y (C_7__0), .A0 (chipmulties_7_cm_nx501), .A1 (
          chipmulties_7_cm_nx503), .A2 (chipmulties_7_cm_nx508), .A3 (
          chipmulties_7_cm_nx518)) ;
    inv01 chipmulties_7_cm_ix502 (.Y (chipmulties_7_cm_nx501), .A (A_7__0)) ;
    oai21 chipmulties_7_cm_ix504 (.Y (chipmulties_7_cm_nx503), .A0 (
          chipmulties_7_cm_nx2), .A1 (A_7__2), .B0 (B_7__0)) ;
    nand02 chipmulties_7_cm_ix3 (.Y (chipmulties_7_cm_nx2), .A0 (
           chipmulties_7_cm_nx506), .A1 (A_7__4)) ;
    inv01 chipmulties_7_cm_ix507 (.Y (chipmulties_7_cm_nx506), .A (A_7__3)) ;
    oai21 chipmulties_7_cm_ix509 (.Y (chipmulties_7_cm_nx508), .A0 (
          chipmulties_7_cm_nx2), .A1 (A_7__1), .B0 (chipmulties_7_cm_nx28)) ;
    aoi21 chipmulties_7_cm_ix29 (.Y (chipmulties_7_cm_nx28), .A0 (
          chipmulties_7_cm_nx511), .A1 (A_7__2), .B0 (chipmulties_7_cm_nx513)) ;
    nand03 chipmulties_7_cm_ix514 (.Y (chipmulties_7_cm_nx513), .A0 (
           chipmulties_7_cm_nx10), .A1 (chipmulties_7_cm_nx12), .A2 (
           chipmulties_7_cm_nx14)) ;
    xnor2 chipmulties_7_cm_ix11 (.Y (chipmulties_7_cm_nx10), .A0 (B_7__3), .A1 (
          B_7__4)) ;
    xnor2 chipmulties_7_cm_ix13 (.Y (chipmulties_7_cm_nx12), .A0 (B_7__2), .A1 (
          B_7__1)) ;
    xnor2 chipmulties_7_cm_ix15 (.Y (chipmulties_7_cm_nx14), .A0 (B_7__3), .A1 (
          B_7__2)) ;
    nor02 chipmulties_7_cm_ix75 (.Y (C_7__1), .A0 (chipmulties_7_cm_nx503), .A1 (
          chipmulties_7_cm_nx523)) ;
    aoi32 chipmulties_7_cm_ix524 (.Y (chipmulties_7_cm_nx523), .A0 (
          chipmulties_7_cm_nx52), .A1 (chipmulties_7_cm_nx54), .A2 (
          chipmulties_7_cm_nx28), .B0 (chipmulties_7_cm_nx46), .B1 (
          chipmulties_7_cm_nx68)) ;
    nor02 chipmulties_7_cm_ix53 (.Y (chipmulties_7_cm_nx52), .A0 (B_7__1), .A1 (
          chipmulties_7_cm_nx46)) ;
    nand02 chipmulties_7_cm_ix47 (.Y (chipmulties_7_cm_nx46), .A0 (A_7__0), .A1 (
           A_7__1)) ;
    nand02 chipmulties_7_cm_ix55 (.Y (chipmulties_7_cm_nx54), .A0 (
           chipmulties_7_cm_nx511), .A1 (chipmulties_7_cm_nx528)) ;
    inv01 chipmulties_7_cm_ix529 (.Y (chipmulties_7_cm_nx528), .A (B_7__4)) ;
    ao32 chipmulties_7_cm_ix69 (.Y (chipmulties_7_cm_nx68), .A0 (B_7__1), .A1 (
         A_7__0), .A2 (chipmulties_7_cm_nx62), .B0 (A_7__1), .B1 (
         chipmulties_7_cm_nx28)) ;
    aoi21 chipmulties_7_cm_ix63 (.Y (chipmulties_7_cm_nx62), .A0 (
          chipmulties_7_cm_nx511), .A1 (chipmulties_7_cm_nx528), .B0 (
          chipmulties_7_cm_nx508)) ;
    nor04 chipmulties_7_cm_ix109 (.Y (C_7__2), .A0 (chipmulties_7_cm_nx508), .A1 (
          chipmulties_7_cm_nx533), .A2 (chipmulties_7_cm_nx535), .A3 (
          chipmulties_7_cm_nx537)) ;
    inv01 chipmulties_7_cm_ix534 (.Y (chipmulties_7_cm_nx533), .A (B_7__0)) ;
    nor03 chipmulties_7_cm_ix536 (.Y (chipmulties_7_cm_nx535), .A0 (A_7__0), .A1 (
          A_7__1), .A2 (A_7__2)) ;
    ao22 chipmulties_7_cm_ix538 (.Y (chipmulties_7_cm_nx537), .A0 (
         chipmulties_7_cm_nx539), .A1 (chipmulties_7_cm_nx543), .B0 (
         chipmulties_7_cm_nx545), .B1 (chipmulties_7_cm_nx547)) ;
    oai21 chipmulties_7_cm_ix540 (.Y (chipmulties_7_cm_nx539), .A0 (A_7__2), .A1 (
          B_7__1), .B0 (chipmulties_7_cm_nx541)) ;
    nor02 chipmulties_7_cm_ix542 (.Y (chipmulties_7_cm_nx541), .A0 (A_7__0), .A1 (
          A_7__1)) ;
    xnor2 chipmulties_7_cm_ix544 (.Y (chipmulties_7_cm_nx543), .A0 (B_7__1), .A1 (
          A_7__2)) ;
    oai22 chipmulties_7_cm_ix546 (.Y (chipmulties_7_cm_nx545), .A0 (
          chipmulties_7_cm_nx2), .A1 (chipmulties_7_cm_nx528), .B0 (
          chipmulties_7_cm_nx506), .B1 (A_7__4)) ;
    nand03 chipmulties_7_cm_ix548 (.Y (chipmulties_7_cm_nx547), .A0 (
           chipmulties_7_cm_nx2), .A1 (B_7__4), .A2 (chipmulties_7_cm_nx46)) ;
    aoi21 chipmulties_7_cm_ix185 (.Y (C_7__3), .A0 (chipmulties_7_cm_nx550), .A1 (
          chipmulties_7_cm_nx569), .B0 (chipmulties_7_cm_nx575)) ;
    oai21 chipmulties_7_cm_ix551 (.Y (chipmulties_7_cm_nx550), .A0 (
          chipmulties_7_cm_nx2), .A1 (A_7__1), .B0 (chipmulties_7_cm_nx178)) ;
    oai22 chipmulties_7_cm_ix179 (.Y (chipmulties_7_cm_nx178), .A0 (
          chipmulties_7_cm_nx553), .A1 (chipmulties_7_cm_nx557), .B0 (
          chipmulties_7_cm_nx528), .B1 (chipmulties_7_cm_nx566)) ;
    aoi21 chipmulties_7_cm_ix554 (.Y (chipmulties_7_cm_nx553), .A0 (
          chipmulties_7_cm_nx555), .A1 (chipmulties_7_cm_nx46), .B0 (A_7__4)) ;
    inv01 chipmulties_7_cm_ix556 (.Y (chipmulties_7_cm_nx555), .A (A_7__2)) ;
    nand02 chipmulties_7_cm_ix558 (.Y (chipmulties_7_cm_nx557), .A0 (
           chipmulties_7_cm_nx528), .A1 (chipmulties_7_cm_nx154)) ;
    oai21 chipmulties_7_cm_ix155 (.Y (chipmulties_7_cm_nx154), .A0 (
          chipmulties_7_cm_nx506), .A1 (A_7__0), .B0 (chipmulties_7_cm_nx560)) ;
    aoi22 chipmulties_7_cm_ix561 (.Y (chipmulties_7_cm_nx560), .A0 (
          chipmulties_7_cm_nx562), .A1 (A_7__3), .B0 (chipmulties_7_cm_nx78), .B1 (
          chipmulties_7_cm_nx130)) ;
    inv01 chipmulties_7_cm_ix563 (.Y (chipmulties_7_cm_nx562), .A (B_7__1)) ;
    aoi32 chipmulties_7_cm_ix567 (.Y (chipmulties_7_cm_nx566), .A0 (
          chipmulties_7_cm_nx164), .A1 (chipmulties_7_cm_nx78), .A2 (
          chipmulties_7_cm_nx130), .B0 (A_7__3), .B1 (chipmulties_7_cm_nx541)) ;
    nand02 chipmulties_7_cm_ix165 (.Y (chipmulties_7_cm_nx164), .A0 (
           chipmulties_7_cm_nx555), .A1 (A_7__4)) ;
    or04 chipmulties_7_cm_ix570 (.Y (chipmulties_7_cm_nx569), .A0 (
         chipmulties_7_cm_nx528), .A1 (A_7__1), .A2 (chipmulties_7_cm_nx560), .A3 (
         chipmulties_7_cm_nx571)) ;
    inv01 chipmulties_7_cm_ix574 (.Y (chipmulties_7_cm_nx573), .A (A_7__4)) ;
    nand03 chipmulties_7_cm_ix576 (.Y (chipmulties_7_cm_nx575), .A0 (
           chipmulties_7_cm_nx118), .A1 (B_7__0), .A2 (chipmulties_7_cm_nx18)) ;
    nand03 chipmulties_7_cm_ix119 (.Y (chipmulties_7_cm_nx118), .A0 (B_7__4), .A1 (
           A_7__2), .A2 (A_7__3)) ;
    nor02 chipmulties_7_cm_ix233 (.Y (C_7__4), .A0 (chipmulties_7_cm_nx575), .A1 (
          chipmulties_7_cm_nx580)) ;
    aoi21 chipmulties_7_cm_ix581 (.Y (chipmulties_7_cm_nx580), .A0 (B_7__1), .A1 (
          chipmulties_7_cm_nx192), .B0 (chipmulties_7_cm_nx228)) ;
    aoi21 chipmulties_7_cm_ix193 (.Y (chipmulties_7_cm_nx192), .A0 (
          chipmulties_7_cm_nx583), .A1 (B_7__4), .B0 (chipmulties_7_cm_nx22)) ;
    oai33 chipmulties_7_cm_ix229 (.Y (chipmulties_7_cm_nx228), .A0 (
          chipmulties_7_cm_nx587), .A1 (chipmulties_7_cm_nx535), .A2 (
          chipmulties_7_cm_nx589), .B0 (B_7__1), .B1 (chipmulties_7_cm_nx573), .B2 (
          chipmulties_7_cm_nx591)) ;
    aoi22 chipmulties_7_cm_ix588 (.Y (chipmulties_7_cm_nx587), .A0 (
          chipmulties_7_cm_nx562), .A1 (chipmulties_7_cm_nx571), .B0 (
          chipmulties_7_cm_nx573), .B1 (chipmulties_7_cm_nx130)) ;
    aoi21 chipmulties_7_cm_ix590 (.Y (chipmulties_7_cm_nx589), .A0 (A_7__2), .A1 (
          A_7__1), .B0 (B_7__4)) ;
    oai21 chipmulties_7_cm_ix592 (.Y (chipmulties_7_cm_nx591), .A0 (
          chipmulties_7_cm_nx46), .A1 (chipmulties_7_cm_nx528), .B0 (A_7__3)) ;
    inv01 chipmulties_7_cm_ix79 (.Y (chipmulties_7_cm_nx78), .A (
          chipmulties_7_cm_nx535)) ;
    inv01 chipmulties_7_cm_ix584 (.Y (chipmulties_7_cm_nx583), .A (
          chipmulties_7_cm_nx46)) ;
    inv01 chipmulties_7_cm_ix23 (.Y (chipmulties_7_cm_nx22), .A (
          chipmulties_7_cm_nx511)) ;
    inv01 chipmulties_7_cm_ix19 (.Y (chipmulties_7_cm_nx18), .A (
          chipmulties_7_cm_nx513)) ;
    inv01 chipmulties_7_cm_ix572 (.Y (chipmulties_7_cm_nx571), .A (
          chipmulties_7_cm_nx2)) ;
    nor02ii chipmulties_7_cm_ix512 (.Y (chipmulties_7_cm_nx511), .A0 (A_7__4), .A1 (
            A_7__3)) ;
    and03 chipmulties_7_cm_ix519 (.Y (chipmulties_7_cm_nx518), .A0 (A_7__3), .A1 (
          chipmulties_7_cm_nx573), .A2 (A_7__1)) ;
    nor02ii chipmulties_7_cm_ix131 (.Y (chipmulties_7_cm_nx130), .A0 (A_7__3), .A1 (
            B_7__1)) ;
    nor04 chipmulties_6_cm_ix41 (.Y (C_6__0), .A0 (chipmulties_6_cm_nx501), .A1 (
          chipmulties_6_cm_nx503), .A2 (chipmulties_6_cm_nx508), .A3 (
          chipmulties_6_cm_nx518)) ;
    inv01 chipmulties_6_cm_ix502 (.Y (chipmulties_6_cm_nx501), .A (A_6__0)) ;
    oai21 chipmulties_6_cm_ix504 (.Y (chipmulties_6_cm_nx503), .A0 (
          chipmulties_6_cm_nx2), .A1 (A_6__2), .B0 (B_6__0)) ;
    nand02 chipmulties_6_cm_ix3 (.Y (chipmulties_6_cm_nx2), .A0 (
           chipmulties_6_cm_nx506), .A1 (A_6__4)) ;
    inv01 chipmulties_6_cm_ix507 (.Y (chipmulties_6_cm_nx506), .A (A_6__3)) ;
    oai21 chipmulties_6_cm_ix509 (.Y (chipmulties_6_cm_nx508), .A0 (
          chipmulties_6_cm_nx2), .A1 (A_6__1), .B0 (chipmulties_6_cm_nx28)) ;
    aoi21 chipmulties_6_cm_ix29 (.Y (chipmulties_6_cm_nx28), .A0 (
          chipmulties_6_cm_nx511), .A1 (A_6__2), .B0 (chipmulties_6_cm_nx513)) ;
    nand03 chipmulties_6_cm_ix514 (.Y (chipmulties_6_cm_nx513), .A0 (
           chipmulties_6_cm_nx10), .A1 (chipmulties_6_cm_nx12), .A2 (
           chipmulties_6_cm_nx14)) ;
    xnor2 chipmulties_6_cm_ix11 (.Y (chipmulties_6_cm_nx10), .A0 (B_6__3), .A1 (
          B_6__4)) ;
    xnor2 chipmulties_6_cm_ix13 (.Y (chipmulties_6_cm_nx12), .A0 (B_6__2), .A1 (
          B_6__1)) ;
    xnor2 chipmulties_6_cm_ix15 (.Y (chipmulties_6_cm_nx14), .A0 (B_6__3), .A1 (
          B_6__2)) ;
    nor02 chipmulties_6_cm_ix75 (.Y (C_6__1), .A0 (chipmulties_6_cm_nx503), .A1 (
          chipmulties_6_cm_nx523)) ;
    aoi32 chipmulties_6_cm_ix524 (.Y (chipmulties_6_cm_nx523), .A0 (
          chipmulties_6_cm_nx52), .A1 (chipmulties_6_cm_nx54), .A2 (
          chipmulties_6_cm_nx28), .B0 (chipmulties_6_cm_nx46), .B1 (
          chipmulties_6_cm_nx68)) ;
    nor02 chipmulties_6_cm_ix53 (.Y (chipmulties_6_cm_nx52), .A0 (B_6__1), .A1 (
          chipmulties_6_cm_nx46)) ;
    nand02 chipmulties_6_cm_ix47 (.Y (chipmulties_6_cm_nx46), .A0 (A_6__0), .A1 (
           A_6__1)) ;
    nand02 chipmulties_6_cm_ix55 (.Y (chipmulties_6_cm_nx54), .A0 (
           chipmulties_6_cm_nx511), .A1 (chipmulties_6_cm_nx528)) ;
    inv01 chipmulties_6_cm_ix529 (.Y (chipmulties_6_cm_nx528), .A (B_6__4)) ;
    ao32 chipmulties_6_cm_ix69 (.Y (chipmulties_6_cm_nx68), .A0 (B_6__1), .A1 (
         A_6__0), .A2 (chipmulties_6_cm_nx62), .B0 (A_6__1), .B1 (
         chipmulties_6_cm_nx28)) ;
    aoi21 chipmulties_6_cm_ix63 (.Y (chipmulties_6_cm_nx62), .A0 (
          chipmulties_6_cm_nx511), .A1 (chipmulties_6_cm_nx528), .B0 (
          chipmulties_6_cm_nx508)) ;
    nor04 chipmulties_6_cm_ix109 (.Y (C_6__2), .A0 (chipmulties_6_cm_nx508), .A1 (
          chipmulties_6_cm_nx533), .A2 (chipmulties_6_cm_nx535), .A3 (
          chipmulties_6_cm_nx537)) ;
    inv01 chipmulties_6_cm_ix534 (.Y (chipmulties_6_cm_nx533), .A (B_6__0)) ;
    nor03 chipmulties_6_cm_ix536 (.Y (chipmulties_6_cm_nx535), .A0 (A_6__0), .A1 (
          A_6__1), .A2 (A_6__2)) ;
    ao22 chipmulties_6_cm_ix538 (.Y (chipmulties_6_cm_nx537), .A0 (
         chipmulties_6_cm_nx539), .A1 (chipmulties_6_cm_nx543), .B0 (
         chipmulties_6_cm_nx545), .B1 (chipmulties_6_cm_nx547)) ;
    oai21 chipmulties_6_cm_ix540 (.Y (chipmulties_6_cm_nx539), .A0 (A_6__2), .A1 (
          B_6__1), .B0 (chipmulties_6_cm_nx541)) ;
    nor02 chipmulties_6_cm_ix542 (.Y (chipmulties_6_cm_nx541), .A0 (A_6__0), .A1 (
          A_6__1)) ;
    xnor2 chipmulties_6_cm_ix544 (.Y (chipmulties_6_cm_nx543), .A0 (B_6__1), .A1 (
          A_6__2)) ;
    oai22 chipmulties_6_cm_ix546 (.Y (chipmulties_6_cm_nx545), .A0 (
          chipmulties_6_cm_nx2), .A1 (chipmulties_6_cm_nx528), .B0 (
          chipmulties_6_cm_nx506), .B1 (A_6__4)) ;
    nand03 chipmulties_6_cm_ix548 (.Y (chipmulties_6_cm_nx547), .A0 (
           chipmulties_6_cm_nx2), .A1 (B_6__4), .A2 (chipmulties_6_cm_nx46)) ;
    aoi21 chipmulties_6_cm_ix185 (.Y (C_6__3), .A0 (chipmulties_6_cm_nx550), .A1 (
          chipmulties_6_cm_nx569), .B0 (chipmulties_6_cm_nx575)) ;
    oai21 chipmulties_6_cm_ix551 (.Y (chipmulties_6_cm_nx550), .A0 (
          chipmulties_6_cm_nx2), .A1 (A_6__1), .B0 (chipmulties_6_cm_nx178)) ;
    oai22 chipmulties_6_cm_ix179 (.Y (chipmulties_6_cm_nx178), .A0 (
          chipmulties_6_cm_nx553), .A1 (chipmulties_6_cm_nx557), .B0 (
          chipmulties_6_cm_nx528), .B1 (chipmulties_6_cm_nx566)) ;
    aoi21 chipmulties_6_cm_ix554 (.Y (chipmulties_6_cm_nx553), .A0 (
          chipmulties_6_cm_nx555), .A1 (chipmulties_6_cm_nx46), .B0 (A_6__4)) ;
    inv01 chipmulties_6_cm_ix556 (.Y (chipmulties_6_cm_nx555), .A (A_6__2)) ;
    nand02 chipmulties_6_cm_ix558 (.Y (chipmulties_6_cm_nx557), .A0 (
           chipmulties_6_cm_nx528), .A1 (chipmulties_6_cm_nx154)) ;
    oai21 chipmulties_6_cm_ix155 (.Y (chipmulties_6_cm_nx154), .A0 (
          chipmulties_6_cm_nx506), .A1 (A_6__0), .B0 (chipmulties_6_cm_nx560)) ;
    aoi22 chipmulties_6_cm_ix561 (.Y (chipmulties_6_cm_nx560), .A0 (
          chipmulties_6_cm_nx562), .A1 (A_6__3), .B0 (chipmulties_6_cm_nx78), .B1 (
          chipmulties_6_cm_nx130)) ;
    inv01 chipmulties_6_cm_ix563 (.Y (chipmulties_6_cm_nx562), .A (B_6__1)) ;
    aoi32 chipmulties_6_cm_ix567 (.Y (chipmulties_6_cm_nx566), .A0 (
          chipmulties_6_cm_nx164), .A1 (chipmulties_6_cm_nx78), .A2 (
          chipmulties_6_cm_nx130), .B0 (A_6__3), .B1 (chipmulties_6_cm_nx541)) ;
    nand02 chipmulties_6_cm_ix165 (.Y (chipmulties_6_cm_nx164), .A0 (
           chipmulties_6_cm_nx555), .A1 (A_6__4)) ;
    or04 chipmulties_6_cm_ix570 (.Y (chipmulties_6_cm_nx569), .A0 (
         chipmulties_6_cm_nx528), .A1 (A_6__1), .A2 (chipmulties_6_cm_nx560), .A3 (
         chipmulties_6_cm_nx571)) ;
    inv01 chipmulties_6_cm_ix574 (.Y (chipmulties_6_cm_nx573), .A (A_6__4)) ;
    nand03 chipmulties_6_cm_ix576 (.Y (chipmulties_6_cm_nx575), .A0 (
           chipmulties_6_cm_nx118), .A1 (B_6__0), .A2 (chipmulties_6_cm_nx18)) ;
    nand03 chipmulties_6_cm_ix119 (.Y (chipmulties_6_cm_nx118), .A0 (B_6__4), .A1 (
           A_6__2), .A2 (A_6__3)) ;
    nor02 chipmulties_6_cm_ix233 (.Y (C_6__4), .A0 (chipmulties_6_cm_nx575), .A1 (
          chipmulties_6_cm_nx580)) ;
    aoi21 chipmulties_6_cm_ix581 (.Y (chipmulties_6_cm_nx580), .A0 (B_6__1), .A1 (
          chipmulties_6_cm_nx192), .B0 (chipmulties_6_cm_nx228)) ;
    aoi21 chipmulties_6_cm_ix193 (.Y (chipmulties_6_cm_nx192), .A0 (
          chipmulties_6_cm_nx583), .A1 (B_6__4), .B0 (chipmulties_6_cm_nx22)) ;
    oai33 chipmulties_6_cm_ix229 (.Y (chipmulties_6_cm_nx228), .A0 (
          chipmulties_6_cm_nx587), .A1 (chipmulties_6_cm_nx535), .A2 (
          chipmulties_6_cm_nx589), .B0 (B_6__1), .B1 (chipmulties_6_cm_nx573), .B2 (
          chipmulties_6_cm_nx591)) ;
    aoi22 chipmulties_6_cm_ix588 (.Y (chipmulties_6_cm_nx587), .A0 (
          chipmulties_6_cm_nx562), .A1 (chipmulties_6_cm_nx571), .B0 (
          chipmulties_6_cm_nx573), .B1 (chipmulties_6_cm_nx130)) ;
    aoi21 chipmulties_6_cm_ix590 (.Y (chipmulties_6_cm_nx589), .A0 (A_6__2), .A1 (
          A_6__1), .B0 (B_6__4)) ;
    oai21 chipmulties_6_cm_ix592 (.Y (chipmulties_6_cm_nx591), .A0 (
          chipmulties_6_cm_nx46), .A1 (chipmulties_6_cm_nx528), .B0 (A_6__3)) ;
    inv01 chipmulties_6_cm_ix79 (.Y (chipmulties_6_cm_nx78), .A (
          chipmulties_6_cm_nx535)) ;
    inv01 chipmulties_6_cm_ix584 (.Y (chipmulties_6_cm_nx583), .A (
          chipmulties_6_cm_nx46)) ;
    inv01 chipmulties_6_cm_ix23 (.Y (chipmulties_6_cm_nx22), .A (
          chipmulties_6_cm_nx511)) ;
    inv01 chipmulties_6_cm_ix19 (.Y (chipmulties_6_cm_nx18), .A (
          chipmulties_6_cm_nx513)) ;
    inv01 chipmulties_6_cm_ix572 (.Y (chipmulties_6_cm_nx571), .A (
          chipmulties_6_cm_nx2)) ;
    nor02ii chipmulties_6_cm_ix512 (.Y (chipmulties_6_cm_nx511), .A0 (A_6__4), .A1 (
            A_6__3)) ;
    and03 chipmulties_6_cm_ix519 (.Y (chipmulties_6_cm_nx518), .A0 (A_6__3), .A1 (
          chipmulties_6_cm_nx573), .A2 (A_6__1)) ;
    nor02ii chipmulties_6_cm_ix131 (.Y (chipmulties_6_cm_nx130), .A0 (A_6__3), .A1 (
            B_6__1)) ;
    nor04 chipmulties_5_cm_ix41 (.Y (C_5__0), .A0 (chipmulties_5_cm_nx501), .A1 (
          chipmulties_5_cm_nx503), .A2 (chipmulties_5_cm_nx508), .A3 (
          chipmulties_5_cm_nx518)) ;
    inv01 chipmulties_5_cm_ix502 (.Y (chipmulties_5_cm_nx501), .A (A_5__0)) ;
    oai21 chipmulties_5_cm_ix504 (.Y (chipmulties_5_cm_nx503), .A0 (
          chipmulties_5_cm_nx2), .A1 (A_5__2), .B0 (B_5__0)) ;
    nand02 chipmulties_5_cm_ix3 (.Y (chipmulties_5_cm_nx2), .A0 (
           chipmulties_5_cm_nx506), .A1 (A_5__4)) ;
    inv01 chipmulties_5_cm_ix507 (.Y (chipmulties_5_cm_nx506), .A (A_5__3)) ;
    oai21 chipmulties_5_cm_ix509 (.Y (chipmulties_5_cm_nx508), .A0 (
          chipmulties_5_cm_nx2), .A1 (A_5__1), .B0 (chipmulties_5_cm_nx28)) ;
    aoi21 chipmulties_5_cm_ix29 (.Y (chipmulties_5_cm_nx28), .A0 (
          chipmulties_5_cm_nx511), .A1 (A_5__2), .B0 (chipmulties_5_cm_nx513)) ;
    nand03 chipmulties_5_cm_ix514 (.Y (chipmulties_5_cm_nx513), .A0 (
           chipmulties_5_cm_nx10), .A1 (chipmulties_5_cm_nx12), .A2 (
           chipmulties_5_cm_nx14)) ;
    xnor2 chipmulties_5_cm_ix11 (.Y (chipmulties_5_cm_nx10), .A0 (B_5__3), .A1 (
          B_5__4)) ;
    xnor2 chipmulties_5_cm_ix13 (.Y (chipmulties_5_cm_nx12), .A0 (B_5__2), .A1 (
          B_5__1)) ;
    xnor2 chipmulties_5_cm_ix15 (.Y (chipmulties_5_cm_nx14), .A0 (B_5__3), .A1 (
          B_5__2)) ;
    nor02 chipmulties_5_cm_ix75 (.Y (C_5__1), .A0 (chipmulties_5_cm_nx503), .A1 (
          chipmulties_5_cm_nx523)) ;
    aoi32 chipmulties_5_cm_ix524 (.Y (chipmulties_5_cm_nx523), .A0 (
          chipmulties_5_cm_nx52), .A1 (chipmulties_5_cm_nx54), .A2 (
          chipmulties_5_cm_nx28), .B0 (chipmulties_5_cm_nx46), .B1 (
          chipmulties_5_cm_nx68)) ;
    nor02 chipmulties_5_cm_ix53 (.Y (chipmulties_5_cm_nx52), .A0 (B_5__1), .A1 (
          chipmulties_5_cm_nx46)) ;
    nand02 chipmulties_5_cm_ix47 (.Y (chipmulties_5_cm_nx46), .A0 (A_5__0), .A1 (
           A_5__1)) ;
    nand02 chipmulties_5_cm_ix55 (.Y (chipmulties_5_cm_nx54), .A0 (
           chipmulties_5_cm_nx511), .A1 (chipmulties_5_cm_nx528)) ;
    inv01 chipmulties_5_cm_ix529 (.Y (chipmulties_5_cm_nx528), .A (B_5__4)) ;
    ao32 chipmulties_5_cm_ix69 (.Y (chipmulties_5_cm_nx68), .A0 (B_5__1), .A1 (
         A_5__0), .A2 (chipmulties_5_cm_nx62), .B0 (A_5__1), .B1 (
         chipmulties_5_cm_nx28)) ;
    aoi21 chipmulties_5_cm_ix63 (.Y (chipmulties_5_cm_nx62), .A0 (
          chipmulties_5_cm_nx511), .A1 (chipmulties_5_cm_nx528), .B0 (
          chipmulties_5_cm_nx508)) ;
    nor04 chipmulties_5_cm_ix109 (.Y (C_5__2), .A0 (chipmulties_5_cm_nx508), .A1 (
          chipmulties_5_cm_nx533), .A2 (chipmulties_5_cm_nx535), .A3 (
          chipmulties_5_cm_nx537)) ;
    inv01 chipmulties_5_cm_ix534 (.Y (chipmulties_5_cm_nx533), .A (B_5__0)) ;
    nor03 chipmulties_5_cm_ix536 (.Y (chipmulties_5_cm_nx535), .A0 (A_5__0), .A1 (
          A_5__1), .A2 (A_5__2)) ;
    ao22 chipmulties_5_cm_ix538 (.Y (chipmulties_5_cm_nx537), .A0 (
         chipmulties_5_cm_nx539), .A1 (chipmulties_5_cm_nx543), .B0 (
         chipmulties_5_cm_nx545), .B1 (chipmulties_5_cm_nx547)) ;
    oai21 chipmulties_5_cm_ix540 (.Y (chipmulties_5_cm_nx539), .A0 (A_5__2), .A1 (
          B_5__1), .B0 (chipmulties_5_cm_nx541)) ;
    nor02 chipmulties_5_cm_ix542 (.Y (chipmulties_5_cm_nx541), .A0 (A_5__0), .A1 (
          A_5__1)) ;
    xnor2 chipmulties_5_cm_ix544 (.Y (chipmulties_5_cm_nx543), .A0 (B_5__1), .A1 (
          A_5__2)) ;
    oai22 chipmulties_5_cm_ix546 (.Y (chipmulties_5_cm_nx545), .A0 (
          chipmulties_5_cm_nx2), .A1 (chipmulties_5_cm_nx528), .B0 (
          chipmulties_5_cm_nx506), .B1 (A_5__4)) ;
    nand03 chipmulties_5_cm_ix548 (.Y (chipmulties_5_cm_nx547), .A0 (
           chipmulties_5_cm_nx2), .A1 (B_5__4), .A2 (chipmulties_5_cm_nx46)) ;
    aoi21 chipmulties_5_cm_ix185 (.Y (C_5__3), .A0 (chipmulties_5_cm_nx550), .A1 (
          chipmulties_5_cm_nx569), .B0 (chipmulties_5_cm_nx575)) ;
    oai21 chipmulties_5_cm_ix551 (.Y (chipmulties_5_cm_nx550), .A0 (
          chipmulties_5_cm_nx2), .A1 (A_5__1), .B0 (chipmulties_5_cm_nx178)) ;
    oai22 chipmulties_5_cm_ix179 (.Y (chipmulties_5_cm_nx178), .A0 (
          chipmulties_5_cm_nx553), .A1 (chipmulties_5_cm_nx557), .B0 (
          chipmulties_5_cm_nx528), .B1 (chipmulties_5_cm_nx566)) ;
    aoi21 chipmulties_5_cm_ix554 (.Y (chipmulties_5_cm_nx553), .A0 (
          chipmulties_5_cm_nx555), .A1 (chipmulties_5_cm_nx46), .B0 (A_5__4)) ;
    inv01 chipmulties_5_cm_ix556 (.Y (chipmulties_5_cm_nx555), .A (A_5__2)) ;
    nand02 chipmulties_5_cm_ix558 (.Y (chipmulties_5_cm_nx557), .A0 (
           chipmulties_5_cm_nx528), .A1 (chipmulties_5_cm_nx154)) ;
    oai21 chipmulties_5_cm_ix155 (.Y (chipmulties_5_cm_nx154), .A0 (
          chipmulties_5_cm_nx506), .A1 (A_5__0), .B0 (chipmulties_5_cm_nx560)) ;
    aoi22 chipmulties_5_cm_ix561 (.Y (chipmulties_5_cm_nx560), .A0 (
          chipmulties_5_cm_nx562), .A1 (A_5__3), .B0 (chipmulties_5_cm_nx78), .B1 (
          chipmulties_5_cm_nx130)) ;
    inv01 chipmulties_5_cm_ix563 (.Y (chipmulties_5_cm_nx562), .A (B_5__1)) ;
    aoi32 chipmulties_5_cm_ix567 (.Y (chipmulties_5_cm_nx566), .A0 (
          chipmulties_5_cm_nx164), .A1 (chipmulties_5_cm_nx78), .A2 (
          chipmulties_5_cm_nx130), .B0 (A_5__3), .B1 (chipmulties_5_cm_nx541)) ;
    nand02 chipmulties_5_cm_ix165 (.Y (chipmulties_5_cm_nx164), .A0 (
           chipmulties_5_cm_nx555), .A1 (A_5__4)) ;
    or04 chipmulties_5_cm_ix570 (.Y (chipmulties_5_cm_nx569), .A0 (
         chipmulties_5_cm_nx528), .A1 (A_5__1), .A2 (chipmulties_5_cm_nx560), .A3 (
         chipmulties_5_cm_nx571)) ;
    inv01 chipmulties_5_cm_ix574 (.Y (chipmulties_5_cm_nx573), .A (A_5__4)) ;
    nand03 chipmulties_5_cm_ix576 (.Y (chipmulties_5_cm_nx575), .A0 (
           chipmulties_5_cm_nx118), .A1 (B_5__0), .A2 (chipmulties_5_cm_nx18)) ;
    nand03 chipmulties_5_cm_ix119 (.Y (chipmulties_5_cm_nx118), .A0 (B_5__4), .A1 (
           A_5__2), .A2 (A_5__3)) ;
    nor02 chipmulties_5_cm_ix233 (.Y (C_5__4), .A0 (chipmulties_5_cm_nx575), .A1 (
          chipmulties_5_cm_nx580)) ;
    aoi21 chipmulties_5_cm_ix581 (.Y (chipmulties_5_cm_nx580), .A0 (B_5__1), .A1 (
          chipmulties_5_cm_nx192), .B0 (chipmulties_5_cm_nx228)) ;
    aoi21 chipmulties_5_cm_ix193 (.Y (chipmulties_5_cm_nx192), .A0 (
          chipmulties_5_cm_nx583), .A1 (B_5__4), .B0 (chipmulties_5_cm_nx22)) ;
    oai33 chipmulties_5_cm_ix229 (.Y (chipmulties_5_cm_nx228), .A0 (
          chipmulties_5_cm_nx587), .A1 (chipmulties_5_cm_nx535), .A2 (
          chipmulties_5_cm_nx589), .B0 (B_5__1), .B1 (chipmulties_5_cm_nx573), .B2 (
          chipmulties_5_cm_nx591)) ;
    aoi22 chipmulties_5_cm_ix588 (.Y (chipmulties_5_cm_nx587), .A0 (
          chipmulties_5_cm_nx562), .A1 (chipmulties_5_cm_nx571), .B0 (
          chipmulties_5_cm_nx573), .B1 (chipmulties_5_cm_nx130)) ;
    aoi21 chipmulties_5_cm_ix590 (.Y (chipmulties_5_cm_nx589), .A0 (A_5__2), .A1 (
          A_5__1), .B0 (B_5__4)) ;
    oai21 chipmulties_5_cm_ix592 (.Y (chipmulties_5_cm_nx591), .A0 (
          chipmulties_5_cm_nx46), .A1 (chipmulties_5_cm_nx528), .B0 (A_5__3)) ;
    inv01 chipmulties_5_cm_ix79 (.Y (chipmulties_5_cm_nx78), .A (
          chipmulties_5_cm_nx535)) ;
    inv01 chipmulties_5_cm_ix584 (.Y (chipmulties_5_cm_nx583), .A (
          chipmulties_5_cm_nx46)) ;
    inv01 chipmulties_5_cm_ix23 (.Y (chipmulties_5_cm_nx22), .A (
          chipmulties_5_cm_nx511)) ;
    inv01 chipmulties_5_cm_ix19 (.Y (chipmulties_5_cm_nx18), .A (
          chipmulties_5_cm_nx513)) ;
    inv01 chipmulties_5_cm_ix572 (.Y (chipmulties_5_cm_nx571), .A (
          chipmulties_5_cm_nx2)) ;
    nor02ii chipmulties_5_cm_ix512 (.Y (chipmulties_5_cm_nx511), .A0 (A_5__4), .A1 (
            A_5__3)) ;
    and03 chipmulties_5_cm_ix519 (.Y (chipmulties_5_cm_nx518), .A0 (A_5__3), .A1 (
          chipmulties_5_cm_nx573), .A2 (A_5__1)) ;
    nor02ii chipmulties_5_cm_ix131 (.Y (chipmulties_5_cm_nx130), .A0 (A_5__3), .A1 (
            B_5__1)) ;
    nor04 chipmulties_4_cm_ix41 (.Y (C_4__0), .A0 (chipmulties_4_cm_nx501), .A1 (
          chipmulties_4_cm_nx503), .A2 (chipmulties_4_cm_nx508), .A3 (
          chipmulties_4_cm_nx518)) ;
    inv01 chipmulties_4_cm_ix502 (.Y (chipmulties_4_cm_nx501), .A (A_4__0)) ;
    oai21 chipmulties_4_cm_ix504 (.Y (chipmulties_4_cm_nx503), .A0 (
          chipmulties_4_cm_nx2), .A1 (A_4__2), .B0 (B_4__0)) ;
    nand02 chipmulties_4_cm_ix3 (.Y (chipmulties_4_cm_nx2), .A0 (
           chipmulties_4_cm_nx506), .A1 (A_4__4)) ;
    inv01 chipmulties_4_cm_ix507 (.Y (chipmulties_4_cm_nx506), .A (A_4__3)) ;
    oai21 chipmulties_4_cm_ix509 (.Y (chipmulties_4_cm_nx508), .A0 (
          chipmulties_4_cm_nx2), .A1 (A_4__1), .B0 (chipmulties_4_cm_nx28)) ;
    aoi21 chipmulties_4_cm_ix29 (.Y (chipmulties_4_cm_nx28), .A0 (
          chipmulties_4_cm_nx511), .A1 (A_4__2), .B0 (chipmulties_4_cm_nx513)) ;
    nand03 chipmulties_4_cm_ix514 (.Y (chipmulties_4_cm_nx513), .A0 (
           chipmulties_4_cm_nx10), .A1 (chipmulties_4_cm_nx12), .A2 (
           chipmulties_4_cm_nx14)) ;
    xnor2 chipmulties_4_cm_ix11 (.Y (chipmulties_4_cm_nx10), .A0 (B_4__3), .A1 (
          B_4__4)) ;
    xnor2 chipmulties_4_cm_ix13 (.Y (chipmulties_4_cm_nx12), .A0 (B_4__2), .A1 (
          B_4__1)) ;
    xnor2 chipmulties_4_cm_ix15 (.Y (chipmulties_4_cm_nx14), .A0 (B_4__3), .A1 (
          B_4__2)) ;
    nor02 chipmulties_4_cm_ix75 (.Y (C_4__1), .A0 (chipmulties_4_cm_nx503), .A1 (
          chipmulties_4_cm_nx523)) ;
    aoi32 chipmulties_4_cm_ix524 (.Y (chipmulties_4_cm_nx523), .A0 (
          chipmulties_4_cm_nx52), .A1 (chipmulties_4_cm_nx54), .A2 (
          chipmulties_4_cm_nx28), .B0 (chipmulties_4_cm_nx46), .B1 (
          chipmulties_4_cm_nx68)) ;
    nor02 chipmulties_4_cm_ix53 (.Y (chipmulties_4_cm_nx52), .A0 (B_4__1), .A1 (
          chipmulties_4_cm_nx46)) ;
    nand02 chipmulties_4_cm_ix47 (.Y (chipmulties_4_cm_nx46), .A0 (A_4__0), .A1 (
           A_4__1)) ;
    nand02 chipmulties_4_cm_ix55 (.Y (chipmulties_4_cm_nx54), .A0 (
           chipmulties_4_cm_nx511), .A1 (chipmulties_4_cm_nx528)) ;
    inv01 chipmulties_4_cm_ix529 (.Y (chipmulties_4_cm_nx528), .A (B_4__4)) ;
    ao32 chipmulties_4_cm_ix69 (.Y (chipmulties_4_cm_nx68), .A0 (B_4__1), .A1 (
         A_4__0), .A2 (chipmulties_4_cm_nx62), .B0 (A_4__1), .B1 (
         chipmulties_4_cm_nx28)) ;
    aoi21 chipmulties_4_cm_ix63 (.Y (chipmulties_4_cm_nx62), .A0 (
          chipmulties_4_cm_nx511), .A1 (chipmulties_4_cm_nx528), .B0 (
          chipmulties_4_cm_nx508)) ;
    nor04 chipmulties_4_cm_ix109 (.Y (C_4__2), .A0 (chipmulties_4_cm_nx508), .A1 (
          chipmulties_4_cm_nx533), .A2 (chipmulties_4_cm_nx535), .A3 (
          chipmulties_4_cm_nx537)) ;
    inv01 chipmulties_4_cm_ix534 (.Y (chipmulties_4_cm_nx533), .A (B_4__0)) ;
    nor03 chipmulties_4_cm_ix536 (.Y (chipmulties_4_cm_nx535), .A0 (A_4__0), .A1 (
          A_4__1), .A2 (A_4__2)) ;
    ao22 chipmulties_4_cm_ix538 (.Y (chipmulties_4_cm_nx537), .A0 (
         chipmulties_4_cm_nx539), .A1 (chipmulties_4_cm_nx543), .B0 (
         chipmulties_4_cm_nx545), .B1 (chipmulties_4_cm_nx547)) ;
    oai21 chipmulties_4_cm_ix540 (.Y (chipmulties_4_cm_nx539), .A0 (A_4__2), .A1 (
          B_4__1), .B0 (chipmulties_4_cm_nx541)) ;
    nor02 chipmulties_4_cm_ix542 (.Y (chipmulties_4_cm_nx541), .A0 (A_4__0), .A1 (
          A_4__1)) ;
    xnor2 chipmulties_4_cm_ix544 (.Y (chipmulties_4_cm_nx543), .A0 (B_4__1), .A1 (
          A_4__2)) ;
    oai22 chipmulties_4_cm_ix546 (.Y (chipmulties_4_cm_nx545), .A0 (
          chipmulties_4_cm_nx2), .A1 (chipmulties_4_cm_nx528), .B0 (
          chipmulties_4_cm_nx506), .B1 (A_4__4)) ;
    nand03 chipmulties_4_cm_ix548 (.Y (chipmulties_4_cm_nx547), .A0 (
           chipmulties_4_cm_nx2), .A1 (B_4__4), .A2 (chipmulties_4_cm_nx46)) ;
    aoi21 chipmulties_4_cm_ix185 (.Y (C_4__3), .A0 (chipmulties_4_cm_nx550), .A1 (
          chipmulties_4_cm_nx569), .B0 (chipmulties_4_cm_nx575)) ;
    oai21 chipmulties_4_cm_ix551 (.Y (chipmulties_4_cm_nx550), .A0 (
          chipmulties_4_cm_nx2), .A1 (A_4__1), .B0 (chipmulties_4_cm_nx178)) ;
    oai22 chipmulties_4_cm_ix179 (.Y (chipmulties_4_cm_nx178), .A0 (
          chipmulties_4_cm_nx553), .A1 (chipmulties_4_cm_nx557), .B0 (
          chipmulties_4_cm_nx528), .B1 (chipmulties_4_cm_nx566)) ;
    aoi21 chipmulties_4_cm_ix554 (.Y (chipmulties_4_cm_nx553), .A0 (
          chipmulties_4_cm_nx555), .A1 (chipmulties_4_cm_nx46), .B0 (A_4__4)) ;
    inv01 chipmulties_4_cm_ix556 (.Y (chipmulties_4_cm_nx555), .A (A_4__2)) ;
    nand02 chipmulties_4_cm_ix558 (.Y (chipmulties_4_cm_nx557), .A0 (
           chipmulties_4_cm_nx528), .A1 (chipmulties_4_cm_nx154)) ;
    oai21 chipmulties_4_cm_ix155 (.Y (chipmulties_4_cm_nx154), .A0 (
          chipmulties_4_cm_nx506), .A1 (A_4__0), .B0 (chipmulties_4_cm_nx560)) ;
    aoi22 chipmulties_4_cm_ix561 (.Y (chipmulties_4_cm_nx560), .A0 (
          chipmulties_4_cm_nx562), .A1 (A_4__3), .B0 (chipmulties_4_cm_nx78), .B1 (
          chipmulties_4_cm_nx130)) ;
    inv01 chipmulties_4_cm_ix563 (.Y (chipmulties_4_cm_nx562), .A (B_4__1)) ;
    aoi32 chipmulties_4_cm_ix567 (.Y (chipmulties_4_cm_nx566), .A0 (
          chipmulties_4_cm_nx164), .A1 (chipmulties_4_cm_nx78), .A2 (
          chipmulties_4_cm_nx130), .B0 (A_4__3), .B1 (chipmulties_4_cm_nx541)) ;
    nand02 chipmulties_4_cm_ix165 (.Y (chipmulties_4_cm_nx164), .A0 (
           chipmulties_4_cm_nx555), .A1 (A_4__4)) ;
    or04 chipmulties_4_cm_ix570 (.Y (chipmulties_4_cm_nx569), .A0 (
         chipmulties_4_cm_nx528), .A1 (A_4__1), .A2 (chipmulties_4_cm_nx560), .A3 (
         chipmulties_4_cm_nx571)) ;
    inv01 chipmulties_4_cm_ix574 (.Y (chipmulties_4_cm_nx573), .A (A_4__4)) ;
    nand03 chipmulties_4_cm_ix576 (.Y (chipmulties_4_cm_nx575), .A0 (
           chipmulties_4_cm_nx118), .A1 (B_4__0), .A2 (chipmulties_4_cm_nx18)) ;
    nand03 chipmulties_4_cm_ix119 (.Y (chipmulties_4_cm_nx118), .A0 (B_4__4), .A1 (
           A_4__2), .A2 (A_4__3)) ;
    nor02 chipmulties_4_cm_ix233 (.Y (C_4__4), .A0 (chipmulties_4_cm_nx575), .A1 (
          chipmulties_4_cm_nx580)) ;
    aoi21 chipmulties_4_cm_ix581 (.Y (chipmulties_4_cm_nx580), .A0 (B_4__1), .A1 (
          chipmulties_4_cm_nx192), .B0 (chipmulties_4_cm_nx228)) ;
    aoi21 chipmulties_4_cm_ix193 (.Y (chipmulties_4_cm_nx192), .A0 (
          chipmulties_4_cm_nx583), .A1 (B_4__4), .B0 (chipmulties_4_cm_nx22)) ;
    oai33 chipmulties_4_cm_ix229 (.Y (chipmulties_4_cm_nx228), .A0 (
          chipmulties_4_cm_nx587), .A1 (chipmulties_4_cm_nx535), .A2 (
          chipmulties_4_cm_nx589), .B0 (B_4__1), .B1 (chipmulties_4_cm_nx573), .B2 (
          chipmulties_4_cm_nx591)) ;
    aoi22 chipmulties_4_cm_ix588 (.Y (chipmulties_4_cm_nx587), .A0 (
          chipmulties_4_cm_nx562), .A1 (chipmulties_4_cm_nx571), .B0 (
          chipmulties_4_cm_nx573), .B1 (chipmulties_4_cm_nx130)) ;
    aoi21 chipmulties_4_cm_ix590 (.Y (chipmulties_4_cm_nx589), .A0 (A_4__2), .A1 (
          A_4__1), .B0 (B_4__4)) ;
    oai21 chipmulties_4_cm_ix592 (.Y (chipmulties_4_cm_nx591), .A0 (
          chipmulties_4_cm_nx46), .A1 (chipmulties_4_cm_nx528), .B0 (A_4__3)) ;
    inv01 chipmulties_4_cm_ix79 (.Y (chipmulties_4_cm_nx78), .A (
          chipmulties_4_cm_nx535)) ;
    inv01 chipmulties_4_cm_ix584 (.Y (chipmulties_4_cm_nx583), .A (
          chipmulties_4_cm_nx46)) ;
    inv01 chipmulties_4_cm_ix23 (.Y (chipmulties_4_cm_nx22), .A (
          chipmulties_4_cm_nx511)) ;
    inv01 chipmulties_4_cm_ix19 (.Y (chipmulties_4_cm_nx18), .A (
          chipmulties_4_cm_nx513)) ;
    inv01 chipmulties_4_cm_ix572 (.Y (chipmulties_4_cm_nx571), .A (
          chipmulties_4_cm_nx2)) ;
    nor02ii chipmulties_4_cm_ix512 (.Y (chipmulties_4_cm_nx511), .A0 (A_4__4), .A1 (
            A_4__3)) ;
    and03 chipmulties_4_cm_ix519 (.Y (chipmulties_4_cm_nx518), .A0 (A_4__3), .A1 (
          chipmulties_4_cm_nx573), .A2 (A_4__1)) ;
    nor02ii chipmulties_4_cm_ix131 (.Y (chipmulties_4_cm_nx130), .A0 (A_4__3), .A1 (
            B_4__1)) ;
    nor04 chipmulties_3_cm_ix41 (.Y (C_3__0), .A0 (chipmulties_3_cm_nx501), .A1 (
          chipmulties_3_cm_nx503), .A2 (chipmulties_3_cm_nx508), .A3 (
          chipmulties_3_cm_nx518)) ;
    inv01 chipmulties_3_cm_ix502 (.Y (chipmulties_3_cm_nx501), .A (A_3__0)) ;
    oai21 chipmulties_3_cm_ix504 (.Y (chipmulties_3_cm_nx503), .A0 (
          chipmulties_3_cm_nx2), .A1 (A_3__2), .B0 (B_3__0)) ;
    nand02 chipmulties_3_cm_ix3 (.Y (chipmulties_3_cm_nx2), .A0 (
           chipmulties_3_cm_nx506), .A1 (A_3__4)) ;
    inv01 chipmulties_3_cm_ix507 (.Y (chipmulties_3_cm_nx506), .A (A_3__3)) ;
    oai21 chipmulties_3_cm_ix509 (.Y (chipmulties_3_cm_nx508), .A0 (
          chipmulties_3_cm_nx2), .A1 (A_3__1), .B0 (chipmulties_3_cm_nx28)) ;
    aoi21 chipmulties_3_cm_ix29 (.Y (chipmulties_3_cm_nx28), .A0 (
          chipmulties_3_cm_nx511), .A1 (A_3__2), .B0 (chipmulties_3_cm_nx513)) ;
    nand03 chipmulties_3_cm_ix514 (.Y (chipmulties_3_cm_nx513), .A0 (
           chipmulties_3_cm_nx10), .A1 (chipmulties_3_cm_nx12), .A2 (
           chipmulties_3_cm_nx14)) ;
    xnor2 chipmulties_3_cm_ix11 (.Y (chipmulties_3_cm_nx10), .A0 (B_3__3), .A1 (
          B_3__4)) ;
    xnor2 chipmulties_3_cm_ix13 (.Y (chipmulties_3_cm_nx12), .A0 (B_3__2), .A1 (
          B_3__1)) ;
    xnor2 chipmulties_3_cm_ix15 (.Y (chipmulties_3_cm_nx14), .A0 (B_3__3), .A1 (
          B_3__2)) ;
    nor02 chipmulties_3_cm_ix75 (.Y (C_3__1), .A0 (chipmulties_3_cm_nx503), .A1 (
          chipmulties_3_cm_nx523)) ;
    aoi32 chipmulties_3_cm_ix524 (.Y (chipmulties_3_cm_nx523), .A0 (
          chipmulties_3_cm_nx52), .A1 (chipmulties_3_cm_nx54), .A2 (
          chipmulties_3_cm_nx28), .B0 (chipmulties_3_cm_nx46), .B1 (
          chipmulties_3_cm_nx68)) ;
    nor02 chipmulties_3_cm_ix53 (.Y (chipmulties_3_cm_nx52), .A0 (B_3__1), .A1 (
          chipmulties_3_cm_nx46)) ;
    nand02 chipmulties_3_cm_ix47 (.Y (chipmulties_3_cm_nx46), .A0 (A_3__0), .A1 (
           A_3__1)) ;
    nand02 chipmulties_3_cm_ix55 (.Y (chipmulties_3_cm_nx54), .A0 (
           chipmulties_3_cm_nx511), .A1 (chipmulties_3_cm_nx528)) ;
    inv01 chipmulties_3_cm_ix529 (.Y (chipmulties_3_cm_nx528), .A (B_3__4)) ;
    ao32 chipmulties_3_cm_ix69 (.Y (chipmulties_3_cm_nx68), .A0 (B_3__1), .A1 (
         A_3__0), .A2 (chipmulties_3_cm_nx62), .B0 (A_3__1), .B1 (
         chipmulties_3_cm_nx28)) ;
    aoi21 chipmulties_3_cm_ix63 (.Y (chipmulties_3_cm_nx62), .A0 (
          chipmulties_3_cm_nx511), .A1 (chipmulties_3_cm_nx528), .B0 (
          chipmulties_3_cm_nx508)) ;
    nor04 chipmulties_3_cm_ix109 (.Y (C_3__2), .A0 (chipmulties_3_cm_nx508), .A1 (
          chipmulties_3_cm_nx533), .A2 (chipmulties_3_cm_nx535), .A3 (
          chipmulties_3_cm_nx537)) ;
    inv01 chipmulties_3_cm_ix534 (.Y (chipmulties_3_cm_nx533), .A (B_3__0)) ;
    nor03 chipmulties_3_cm_ix536 (.Y (chipmulties_3_cm_nx535), .A0 (A_3__0), .A1 (
          A_3__1), .A2 (A_3__2)) ;
    ao22 chipmulties_3_cm_ix538 (.Y (chipmulties_3_cm_nx537), .A0 (
         chipmulties_3_cm_nx539), .A1 (chipmulties_3_cm_nx543), .B0 (
         chipmulties_3_cm_nx545), .B1 (chipmulties_3_cm_nx547)) ;
    oai21 chipmulties_3_cm_ix540 (.Y (chipmulties_3_cm_nx539), .A0 (A_3__2), .A1 (
          B_3__1), .B0 (chipmulties_3_cm_nx541)) ;
    nor02 chipmulties_3_cm_ix542 (.Y (chipmulties_3_cm_nx541), .A0 (A_3__0), .A1 (
          A_3__1)) ;
    xnor2 chipmulties_3_cm_ix544 (.Y (chipmulties_3_cm_nx543), .A0 (B_3__1), .A1 (
          A_3__2)) ;
    oai22 chipmulties_3_cm_ix546 (.Y (chipmulties_3_cm_nx545), .A0 (
          chipmulties_3_cm_nx2), .A1 (chipmulties_3_cm_nx528), .B0 (
          chipmulties_3_cm_nx506), .B1 (A_3__4)) ;
    nand03 chipmulties_3_cm_ix548 (.Y (chipmulties_3_cm_nx547), .A0 (
           chipmulties_3_cm_nx2), .A1 (B_3__4), .A2 (chipmulties_3_cm_nx46)) ;
    aoi21 chipmulties_3_cm_ix185 (.Y (C_3__3), .A0 (chipmulties_3_cm_nx550), .A1 (
          chipmulties_3_cm_nx569), .B0 (chipmulties_3_cm_nx575)) ;
    oai21 chipmulties_3_cm_ix551 (.Y (chipmulties_3_cm_nx550), .A0 (
          chipmulties_3_cm_nx2), .A1 (A_3__1), .B0 (chipmulties_3_cm_nx178)) ;
    oai22 chipmulties_3_cm_ix179 (.Y (chipmulties_3_cm_nx178), .A0 (
          chipmulties_3_cm_nx553), .A1 (chipmulties_3_cm_nx557), .B0 (
          chipmulties_3_cm_nx528), .B1 (chipmulties_3_cm_nx566)) ;
    aoi21 chipmulties_3_cm_ix554 (.Y (chipmulties_3_cm_nx553), .A0 (
          chipmulties_3_cm_nx555), .A1 (chipmulties_3_cm_nx46), .B0 (A_3__4)) ;
    inv01 chipmulties_3_cm_ix556 (.Y (chipmulties_3_cm_nx555), .A (A_3__2)) ;
    nand02 chipmulties_3_cm_ix558 (.Y (chipmulties_3_cm_nx557), .A0 (
           chipmulties_3_cm_nx528), .A1 (chipmulties_3_cm_nx154)) ;
    oai21 chipmulties_3_cm_ix155 (.Y (chipmulties_3_cm_nx154), .A0 (
          chipmulties_3_cm_nx506), .A1 (A_3__0), .B0 (chipmulties_3_cm_nx560)) ;
    aoi22 chipmulties_3_cm_ix561 (.Y (chipmulties_3_cm_nx560), .A0 (
          chipmulties_3_cm_nx562), .A1 (A_3__3), .B0 (chipmulties_3_cm_nx78), .B1 (
          chipmulties_3_cm_nx130)) ;
    inv01 chipmulties_3_cm_ix563 (.Y (chipmulties_3_cm_nx562), .A (B_3__1)) ;
    aoi32 chipmulties_3_cm_ix567 (.Y (chipmulties_3_cm_nx566), .A0 (
          chipmulties_3_cm_nx164), .A1 (chipmulties_3_cm_nx78), .A2 (
          chipmulties_3_cm_nx130), .B0 (A_3__3), .B1 (chipmulties_3_cm_nx541)) ;
    nand02 chipmulties_3_cm_ix165 (.Y (chipmulties_3_cm_nx164), .A0 (
           chipmulties_3_cm_nx555), .A1 (A_3__4)) ;
    or04 chipmulties_3_cm_ix570 (.Y (chipmulties_3_cm_nx569), .A0 (
         chipmulties_3_cm_nx528), .A1 (A_3__1), .A2 (chipmulties_3_cm_nx560), .A3 (
         chipmulties_3_cm_nx571)) ;
    inv01 chipmulties_3_cm_ix574 (.Y (chipmulties_3_cm_nx573), .A (A_3__4)) ;
    nand03 chipmulties_3_cm_ix576 (.Y (chipmulties_3_cm_nx575), .A0 (
           chipmulties_3_cm_nx118), .A1 (B_3__0), .A2 (chipmulties_3_cm_nx18)) ;
    nand03 chipmulties_3_cm_ix119 (.Y (chipmulties_3_cm_nx118), .A0 (B_3__4), .A1 (
           A_3__2), .A2 (A_3__3)) ;
    nor02 chipmulties_3_cm_ix233 (.Y (C_3__4), .A0 (chipmulties_3_cm_nx575), .A1 (
          chipmulties_3_cm_nx580)) ;
    aoi21 chipmulties_3_cm_ix581 (.Y (chipmulties_3_cm_nx580), .A0 (B_3__1), .A1 (
          chipmulties_3_cm_nx192), .B0 (chipmulties_3_cm_nx228)) ;
    aoi21 chipmulties_3_cm_ix193 (.Y (chipmulties_3_cm_nx192), .A0 (
          chipmulties_3_cm_nx583), .A1 (B_3__4), .B0 (chipmulties_3_cm_nx22)) ;
    oai33 chipmulties_3_cm_ix229 (.Y (chipmulties_3_cm_nx228), .A0 (
          chipmulties_3_cm_nx587), .A1 (chipmulties_3_cm_nx535), .A2 (
          chipmulties_3_cm_nx589), .B0 (B_3__1), .B1 (chipmulties_3_cm_nx573), .B2 (
          chipmulties_3_cm_nx591)) ;
    aoi22 chipmulties_3_cm_ix588 (.Y (chipmulties_3_cm_nx587), .A0 (
          chipmulties_3_cm_nx562), .A1 (chipmulties_3_cm_nx571), .B0 (
          chipmulties_3_cm_nx573), .B1 (chipmulties_3_cm_nx130)) ;
    aoi21 chipmulties_3_cm_ix590 (.Y (chipmulties_3_cm_nx589), .A0 (A_3__2), .A1 (
          A_3__1), .B0 (B_3__4)) ;
    oai21 chipmulties_3_cm_ix592 (.Y (chipmulties_3_cm_nx591), .A0 (
          chipmulties_3_cm_nx46), .A1 (chipmulties_3_cm_nx528), .B0 (A_3__3)) ;
    inv01 chipmulties_3_cm_ix79 (.Y (chipmulties_3_cm_nx78), .A (
          chipmulties_3_cm_nx535)) ;
    inv01 chipmulties_3_cm_ix584 (.Y (chipmulties_3_cm_nx583), .A (
          chipmulties_3_cm_nx46)) ;
    inv01 chipmulties_3_cm_ix23 (.Y (chipmulties_3_cm_nx22), .A (
          chipmulties_3_cm_nx511)) ;
    inv01 chipmulties_3_cm_ix19 (.Y (chipmulties_3_cm_nx18), .A (
          chipmulties_3_cm_nx513)) ;
    inv01 chipmulties_3_cm_ix572 (.Y (chipmulties_3_cm_nx571), .A (
          chipmulties_3_cm_nx2)) ;
    nor02ii chipmulties_3_cm_ix512 (.Y (chipmulties_3_cm_nx511), .A0 (A_3__4), .A1 (
            A_3__3)) ;
    and03 chipmulties_3_cm_ix519 (.Y (chipmulties_3_cm_nx518), .A0 (A_3__3), .A1 (
          chipmulties_3_cm_nx573), .A2 (A_3__1)) ;
    nor02ii chipmulties_3_cm_ix131 (.Y (chipmulties_3_cm_nx130), .A0 (A_3__3), .A1 (
            B_3__1)) ;
    nor04 chipmulties_2_cm_ix41 (.Y (C_2__0), .A0 (chipmulties_2_cm_nx501), .A1 (
          chipmulties_2_cm_nx503), .A2 (chipmulties_2_cm_nx508), .A3 (
          chipmulties_2_cm_nx518)) ;
    inv01 chipmulties_2_cm_ix502 (.Y (chipmulties_2_cm_nx501), .A (A_2__0)) ;
    oai21 chipmulties_2_cm_ix504 (.Y (chipmulties_2_cm_nx503), .A0 (
          chipmulties_2_cm_nx2), .A1 (A_2__2), .B0 (B_2__0)) ;
    nand02 chipmulties_2_cm_ix3 (.Y (chipmulties_2_cm_nx2), .A0 (
           chipmulties_2_cm_nx506), .A1 (A_2__4)) ;
    inv01 chipmulties_2_cm_ix507 (.Y (chipmulties_2_cm_nx506), .A (A_2__3)) ;
    oai21 chipmulties_2_cm_ix509 (.Y (chipmulties_2_cm_nx508), .A0 (
          chipmulties_2_cm_nx2), .A1 (A_2__1), .B0 (chipmulties_2_cm_nx28)) ;
    aoi21 chipmulties_2_cm_ix29 (.Y (chipmulties_2_cm_nx28), .A0 (
          chipmulties_2_cm_nx511), .A1 (A_2__2), .B0 (chipmulties_2_cm_nx513)) ;
    nand03 chipmulties_2_cm_ix514 (.Y (chipmulties_2_cm_nx513), .A0 (
           chipmulties_2_cm_nx10), .A1 (chipmulties_2_cm_nx12), .A2 (
           chipmulties_2_cm_nx14)) ;
    xnor2 chipmulties_2_cm_ix11 (.Y (chipmulties_2_cm_nx10), .A0 (B_2__3), .A1 (
          B_2__4)) ;
    xnor2 chipmulties_2_cm_ix13 (.Y (chipmulties_2_cm_nx12), .A0 (B_2__2), .A1 (
          B_2__1)) ;
    xnor2 chipmulties_2_cm_ix15 (.Y (chipmulties_2_cm_nx14), .A0 (B_2__3), .A1 (
          B_2__2)) ;
    nor02 chipmulties_2_cm_ix75 (.Y (C_2__1), .A0 (chipmulties_2_cm_nx503), .A1 (
          chipmulties_2_cm_nx523)) ;
    aoi32 chipmulties_2_cm_ix524 (.Y (chipmulties_2_cm_nx523), .A0 (
          chipmulties_2_cm_nx52), .A1 (chipmulties_2_cm_nx54), .A2 (
          chipmulties_2_cm_nx28), .B0 (chipmulties_2_cm_nx46), .B1 (
          chipmulties_2_cm_nx68)) ;
    nor02 chipmulties_2_cm_ix53 (.Y (chipmulties_2_cm_nx52), .A0 (B_2__1), .A1 (
          chipmulties_2_cm_nx46)) ;
    nand02 chipmulties_2_cm_ix47 (.Y (chipmulties_2_cm_nx46), .A0 (A_2__0), .A1 (
           A_2__1)) ;
    nand02 chipmulties_2_cm_ix55 (.Y (chipmulties_2_cm_nx54), .A0 (
           chipmulties_2_cm_nx511), .A1 (chipmulties_2_cm_nx528)) ;
    inv01 chipmulties_2_cm_ix529 (.Y (chipmulties_2_cm_nx528), .A (B_2__4)) ;
    ao32 chipmulties_2_cm_ix69 (.Y (chipmulties_2_cm_nx68), .A0 (B_2__1), .A1 (
         A_2__0), .A2 (chipmulties_2_cm_nx62), .B0 (A_2__1), .B1 (
         chipmulties_2_cm_nx28)) ;
    aoi21 chipmulties_2_cm_ix63 (.Y (chipmulties_2_cm_nx62), .A0 (
          chipmulties_2_cm_nx511), .A1 (chipmulties_2_cm_nx528), .B0 (
          chipmulties_2_cm_nx508)) ;
    nor04 chipmulties_2_cm_ix109 (.Y (C_2__2), .A0 (chipmulties_2_cm_nx508), .A1 (
          chipmulties_2_cm_nx533), .A2 (chipmulties_2_cm_nx535), .A3 (
          chipmulties_2_cm_nx537)) ;
    inv01 chipmulties_2_cm_ix534 (.Y (chipmulties_2_cm_nx533), .A (B_2__0)) ;
    nor03 chipmulties_2_cm_ix536 (.Y (chipmulties_2_cm_nx535), .A0 (A_2__0), .A1 (
          A_2__1), .A2 (A_2__2)) ;
    ao22 chipmulties_2_cm_ix538 (.Y (chipmulties_2_cm_nx537), .A0 (
         chipmulties_2_cm_nx539), .A1 (chipmulties_2_cm_nx543), .B0 (
         chipmulties_2_cm_nx545), .B1 (chipmulties_2_cm_nx547)) ;
    oai21 chipmulties_2_cm_ix540 (.Y (chipmulties_2_cm_nx539), .A0 (A_2__2), .A1 (
          B_2__1), .B0 (chipmulties_2_cm_nx541)) ;
    nor02 chipmulties_2_cm_ix542 (.Y (chipmulties_2_cm_nx541), .A0 (A_2__0), .A1 (
          A_2__1)) ;
    xnor2 chipmulties_2_cm_ix544 (.Y (chipmulties_2_cm_nx543), .A0 (B_2__1), .A1 (
          A_2__2)) ;
    oai22 chipmulties_2_cm_ix546 (.Y (chipmulties_2_cm_nx545), .A0 (
          chipmulties_2_cm_nx2), .A1 (chipmulties_2_cm_nx528), .B0 (
          chipmulties_2_cm_nx506), .B1 (A_2__4)) ;
    nand03 chipmulties_2_cm_ix548 (.Y (chipmulties_2_cm_nx547), .A0 (
           chipmulties_2_cm_nx2), .A1 (B_2__4), .A2 (chipmulties_2_cm_nx46)) ;
    aoi21 chipmulties_2_cm_ix185 (.Y (C_2__3), .A0 (chipmulties_2_cm_nx550), .A1 (
          chipmulties_2_cm_nx569), .B0 (chipmulties_2_cm_nx575)) ;
    oai21 chipmulties_2_cm_ix551 (.Y (chipmulties_2_cm_nx550), .A0 (
          chipmulties_2_cm_nx2), .A1 (A_2__1), .B0 (chipmulties_2_cm_nx178)) ;
    oai22 chipmulties_2_cm_ix179 (.Y (chipmulties_2_cm_nx178), .A0 (
          chipmulties_2_cm_nx553), .A1 (chipmulties_2_cm_nx557), .B0 (
          chipmulties_2_cm_nx528), .B1 (chipmulties_2_cm_nx566)) ;
    aoi21 chipmulties_2_cm_ix554 (.Y (chipmulties_2_cm_nx553), .A0 (
          chipmulties_2_cm_nx555), .A1 (chipmulties_2_cm_nx46), .B0 (A_2__4)) ;
    inv01 chipmulties_2_cm_ix556 (.Y (chipmulties_2_cm_nx555), .A (A_2__2)) ;
    nand02 chipmulties_2_cm_ix558 (.Y (chipmulties_2_cm_nx557), .A0 (
           chipmulties_2_cm_nx528), .A1 (chipmulties_2_cm_nx154)) ;
    oai21 chipmulties_2_cm_ix155 (.Y (chipmulties_2_cm_nx154), .A0 (
          chipmulties_2_cm_nx506), .A1 (A_2__0), .B0 (chipmulties_2_cm_nx560)) ;
    aoi22 chipmulties_2_cm_ix561 (.Y (chipmulties_2_cm_nx560), .A0 (
          chipmulties_2_cm_nx562), .A1 (A_2__3), .B0 (chipmulties_2_cm_nx78), .B1 (
          chipmulties_2_cm_nx130)) ;
    inv01 chipmulties_2_cm_ix563 (.Y (chipmulties_2_cm_nx562), .A (B_2__1)) ;
    aoi32 chipmulties_2_cm_ix567 (.Y (chipmulties_2_cm_nx566), .A0 (
          chipmulties_2_cm_nx164), .A1 (chipmulties_2_cm_nx78), .A2 (
          chipmulties_2_cm_nx130), .B0 (A_2__3), .B1 (chipmulties_2_cm_nx541)) ;
    nand02 chipmulties_2_cm_ix165 (.Y (chipmulties_2_cm_nx164), .A0 (
           chipmulties_2_cm_nx555), .A1 (A_2__4)) ;
    or04 chipmulties_2_cm_ix570 (.Y (chipmulties_2_cm_nx569), .A0 (
         chipmulties_2_cm_nx528), .A1 (A_2__1), .A2 (chipmulties_2_cm_nx560), .A3 (
         chipmulties_2_cm_nx571)) ;
    inv01 chipmulties_2_cm_ix574 (.Y (chipmulties_2_cm_nx573), .A (A_2__4)) ;
    nand03 chipmulties_2_cm_ix576 (.Y (chipmulties_2_cm_nx575), .A0 (
           chipmulties_2_cm_nx118), .A1 (B_2__0), .A2 (chipmulties_2_cm_nx18)) ;
    nand03 chipmulties_2_cm_ix119 (.Y (chipmulties_2_cm_nx118), .A0 (B_2__4), .A1 (
           A_2__2), .A2 (A_2__3)) ;
    nor02 chipmulties_2_cm_ix233 (.Y (C_2__4), .A0 (chipmulties_2_cm_nx575), .A1 (
          chipmulties_2_cm_nx580)) ;
    aoi21 chipmulties_2_cm_ix581 (.Y (chipmulties_2_cm_nx580), .A0 (B_2__1), .A1 (
          chipmulties_2_cm_nx192), .B0 (chipmulties_2_cm_nx228)) ;
    aoi21 chipmulties_2_cm_ix193 (.Y (chipmulties_2_cm_nx192), .A0 (
          chipmulties_2_cm_nx583), .A1 (B_2__4), .B0 (chipmulties_2_cm_nx22)) ;
    oai33 chipmulties_2_cm_ix229 (.Y (chipmulties_2_cm_nx228), .A0 (
          chipmulties_2_cm_nx587), .A1 (chipmulties_2_cm_nx535), .A2 (
          chipmulties_2_cm_nx589), .B0 (B_2__1), .B1 (chipmulties_2_cm_nx573), .B2 (
          chipmulties_2_cm_nx591)) ;
    aoi22 chipmulties_2_cm_ix588 (.Y (chipmulties_2_cm_nx587), .A0 (
          chipmulties_2_cm_nx562), .A1 (chipmulties_2_cm_nx571), .B0 (
          chipmulties_2_cm_nx573), .B1 (chipmulties_2_cm_nx130)) ;
    aoi21 chipmulties_2_cm_ix590 (.Y (chipmulties_2_cm_nx589), .A0 (A_2__2), .A1 (
          A_2__1), .B0 (B_2__4)) ;
    oai21 chipmulties_2_cm_ix592 (.Y (chipmulties_2_cm_nx591), .A0 (
          chipmulties_2_cm_nx46), .A1 (chipmulties_2_cm_nx528), .B0 (A_2__3)) ;
    inv01 chipmulties_2_cm_ix79 (.Y (chipmulties_2_cm_nx78), .A (
          chipmulties_2_cm_nx535)) ;
    inv01 chipmulties_2_cm_ix584 (.Y (chipmulties_2_cm_nx583), .A (
          chipmulties_2_cm_nx46)) ;
    inv01 chipmulties_2_cm_ix23 (.Y (chipmulties_2_cm_nx22), .A (
          chipmulties_2_cm_nx511)) ;
    inv01 chipmulties_2_cm_ix19 (.Y (chipmulties_2_cm_nx18), .A (
          chipmulties_2_cm_nx513)) ;
    inv01 chipmulties_2_cm_ix572 (.Y (chipmulties_2_cm_nx571), .A (
          chipmulties_2_cm_nx2)) ;
    nor02ii chipmulties_2_cm_ix512 (.Y (chipmulties_2_cm_nx511), .A0 (A_2__4), .A1 (
            A_2__3)) ;
    and03 chipmulties_2_cm_ix519 (.Y (chipmulties_2_cm_nx518), .A0 (A_2__3), .A1 (
          chipmulties_2_cm_nx573), .A2 (A_2__1)) ;
    nor02ii chipmulties_2_cm_ix131 (.Y (chipmulties_2_cm_nx130), .A0 (A_2__3), .A1 (
            B_2__1)) ;
    nor04 chipmulties_1_cm_ix41 (.Y (C_1__0), .A0 (chipmulties_1_cm_nx501), .A1 (
          chipmulties_1_cm_nx503), .A2 (chipmulties_1_cm_nx508), .A3 (
          chipmulties_1_cm_nx518)) ;
    inv01 chipmulties_1_cm_ix502 (.Y (chipmulties_1_cm_nx501), .A (A_1__0)) ;
    oai21 chipmulties_1_cm_ix504 (.Y (chipmulties_1_cm_nx503), .A0 (
          chipmulties_1_cm_nx2), .A1 (A_1__2), .B0 (B_1__0)) ;
    nand02 chipmulties_1_cm_ix3 (.Y (chipmulties_1_cm_nx2), .A0 (
           chipmulties_1_cm_nx506), .A1 (A_1__4)) ;
    inv01 chipmulties_1_cm_ix507 (.Y (chipmulties_1_cm_nx506), .A (A_1__3)) ;
    oai21 chipmulties_1_cm_ix509 (.Y (chipmulties_1_cm_nx508), .A0 (
          chipmulties_1_cm_nx2), .A1 (A_1__1), .B0 (chipmulties_1_cm_nx28)) ;
    aoi21 chipmulties_1_cm_ix29 (.Y (chipmulties_1_cm_nx28), .A0 (
          chipmulties_1_cm_nx511), .A1 (A_1__2), .B0 (chipmulties_1_cm_nx513)) ;
    nand03 chipmulties_1_cm_ix514 (.Y (chipmulties_1_cm_nx513), .A0 (
           chipmulties_1_cm_nx10), .A1 (chipmulties_1_cm_nx12), .A2 (
           chipmulties_1_cm_nx14)) ;
    xnor2 chipmulties_1_cm_ix11 (.Y (chipmulties_1_cm_nx10), .A0 (B_1__3), .A1 (
          B_1__4)) ;
    xnor2 chipmulties_1_cm_ix13 (.Y (chipmulties_1_cm_nx12), .A0 (B_1__2), .A1 (
          B_1__1)) ;
    xnor2 chipmulties_1_cm_ix15 (.Y (chipmulties_1_cm_nx14), .A0 (B_1__3), .A1 (
          B_1__2)) ;
    nor02 chipmulties_1_cm_ix75 (.Y (C_1__1), .A0 (chipmulties_1_cm_nx503), .A1 (
          chipmulties_1_cm_nx523)) ;
    aoi32 chipmulties_1_cm_ix524 (.Y (chipmulties_1_cm_nx523), .A0 (
          chipmulties_1_cm_nx52), .A1 (chipmulties_1_cm_nx54), .A2 (
          chipmulties_1_cm_nx28), .B0 (chipmulties_1_cm_nx46), .B1 (
          chipmulties_1_cm_nx68)) ;
    nor02 chipmulties_1_cm_ix53 (.Y (chipmulties_1_cm_nx52), .A0 (B_1__1), .A1 (
          chipmulties_1_cm_nx46)) ;
    nand02 chipmulties_1_cm_ix47 (.Y (chipmulties_1_cm_nx46), .A0 (A_1__0), .A1 (
           A_1__1)) ;
    nand02 chipmulties_1_cm_ix55 (.Y (chipmulties_1_cm_nx54), .A0 (
           chipmulties_1_cm_nx511), .A1 (chipmulties_1_cm_nx528)) ;
    inv01 chipmulties_1_cm_ix529 (.Y (chipmulties_1_cm_nx528), .A (B_1__4)) ;
    ao32 chipmulties_1_cm_ix69 (.Y (chipmulties_1_cm_nx68), .A0 (B_1__1), .A1 (
         A_1__0), .A2 (chipmulties_1_cm_nx62), .B0 (A_1__1), .B1 (
         chipmulties_1_cm_nx28)) ;
    aoi21 chipmulties_1_cm_ix63 (.Y (chipmulties_1_cm_nx62), .A0 (
          chipmulties_1_cm_nx511), .A1 (chipmulties_1_cm_nx528), .B0 (
          chipmulties_1_cm_nx508)) ;
    nor04 chipmulties_1_cm_ix109 (.Y (C_1__2), .A0 (chipmulties_1_cm_nx508), .A1 (
          chipmulties_1_cm_nx533), .A2 (chipmulties_1_cm_nx535), .A3 (
          chipmulties_1_cm_nx537)) ;
    inv01 chipmulties_1_cm_ix534 (.Y (chipmulties_1_cm_nx533), .A (B_1__0)) ;
    nor03 chipmulties_1_cm_ix536 (.Y (chipmulties_1_cm_nx535), .A0 (A_1__0), .A1 (
          A_1__1), .A2 (A_1__2)) ;
    ao22 chipmulties_1_cm_ix538 (.Y (chipmulties_1_cm_nx537), .A0 (
         chipmulties_1_cm_nx539), .A1 (chipmulties_1_cm_nx543), .B0 (
         chipmulties_1_cm_nx545), .B1 (chipmulties_1_cm_nx547)) ;
    oai21 chipmulties_1_cm_ix540 (.Y (chipmulties_1_cm_nx539), .A0 (A_1__2), .A1 (
          B_1__1), .B0 (chipmulties_1_cm_nx541)) ;
    nor02 chipmulties_1_cm_ix542 (.Y (chipmulties_1_cm_nx541), .A0 (A_1__0), .A1 (
          A_1__1)) ;
    xnor2 chipmulties_1_cm_ix544 (.Y (chipmulties_1_cm_nx543), .A0 (B_1__1), .A1 (
          A_1__2)) ;
    oai22 chipmulties_1_cm_ix546 (.Y (chipmulties_1_cm_nx545), .A0 (
          chipmulties_1_cm_nx2), .A1 (chipmulties_1_cm_nx528), .B0 (
          chipmulties_1_cm_nx506), .B1 (A_1__4)) ;
    nand03 chipmulties_1_cm_ix548 (.Y (chipmulties_1_cm_nx547), .A0 (
           chipmulties_1_cm_nx2), .A1 (B_1__4), .A2 (chipmulties_1_cm_nx46)) ;
    aoi21 chipmulties_1_cm_ix185 (.Y (C_1__3), .A0 (chipmulties_1_cm_nx550), .A1 (
          chipmulties_1_cm_nx569), .B0 (chipmulties_1_cm_nx575)) ;
    oai21 chipmulties_1_cm_ix551 (.Y (chipmulties_1_cm_nx550), .A0 (
          chipmulties_1_cm_nx2), .A1 (A_1__1), .B0 (chipmulties_1_cm_nx178)) ;
    oai22 chipmulties_1_cm_ix179 (.Y (chipmulties_1_cm_nx178), .A0 (
          chipmulties_1_cm_nx553), .A1 (chipmulties_1_cm_nx557), .B0 (
          chipmulties_1_cm_nx528), .B1 (chipmulties_1_cm_nx566)) ;
    aoi21 chipmulties_1_cm_ix554 (.Y (chipmulties_1_cm_nx553), .A0 (
          chipmulties_1_cm_nx555), .A1 (chipmulties_1_cm_nx46), .B0 (A_1__4)) ;
    inv01 chipmulties_1_cm_ix556 (.Y (chipmulties_1_cm_nx555), .A (A_1__2)) ;
    nand02 chipmulties_1_cm_ix558 (.Y (chipmulties_1_cm_nx557), .A0 (
           chipmulties_1_cm_nx528), .A1 (chipmulties_1_cm_nx154)) ;
    oai21 chipmulties_1_cm_ix155 (.Y (chipmulties_1_cm_nx154), .A0 (
          chipmulties_1_cm_nx506), .A1 (A_1__0), .B0 (chipmulties_1_cm_nx560)) ;
    aoi22 chipmulties_1_cm_ix561 (.Y (chipmulties_1_cm_nx560), .A0 (
          chipmulties_1_cm_nx562), .A1 (A_1__3), .B0 (chipmulties_1_cm_nx78), .B1 (
          chipmulties_1_cm_nx130)) ;
    inv01 chipmulties_1_cm_ix563 (.Y (chipmulties_1_cm_nx562), .A (B_1__1)) ;
    aoi32 chipmulties_1_cm_ix567 (.Y (chipmulties_1_cm_nx566), .A0 (
          chipmulties_1_cm_nx164), .A1 (chipmulties_1_cm_nx78), .A2 (
          chipmulties_1_cm_nx130), .B0 (A_1__3), .B1 (chipmulties_1_cm_nx541)) ;
    nand02 chipmulties_1_cm_ix165 (.Y (chipmulties_1_cm_nx164), .A0 (
           chipmulties_1_cm_nx555), .A1 (A_1__4)) ;
    or04 chipmulties_1_cm_ix570 (.Y (chipmulties_1_cm_nx569), .A0 (
         chipmulties_1_cm_nx528), .A1 (A_1__1), .A2 (chipmulties_1_cm_nx560), .A3 (
         chipmulties_1_cm_nx571)) ;
    inv01 chipmulties_1_cm_ix574 (.Y (chipmulties_1_cm_nx573), .A (A_1__4)) ;
    nand03 chipmulties_1_cm_ix576 (.Y (chipmulties_1_cm_nx575), .A0 (
           chipmulties_1_cm_nx118), .A1 (B_1__0), .A2 (chipmulties_1_cm_nx18)) ;
    nand03 chipmulties_1_cm_ix119 (.Y (chipmulties_1_cm_nx118), .A0 (B_1__4), .A1 (
           A_1__2), .A2 (A_1__3)) ;
    nor02 chipmulties_1_cm_ix233 (.Y (C_1__4), .A0 (chipmulties_1_cm_nx575), .A1 (
          chipmulties_1_cm_nx580)) ;
    aoi21 chipmulties_1_cm_ix581 (.Y (chipmulties_1_cm_nx580), .A0 (B_1__1), .A1 (
          chipmulties_1_cm_nx192), .B0 (chipmulties_1_cm_nx228)) ;
    aoi21 chipmulties_1_cm_ix193 (.Y (chipmulties_1_cm_nx192), .A0 (
          chipmulties_1_cm_nx583), .A1 (B_1__4), .B0 (chipmulties_1_cm_nx22)) ;
    oai33 chipmulties_1_cm_ix229 (.Y (chipmulties_1_cm_nx228), .A0 (
          chipmulties_1_cm_nx587), .A1 (chipmulties_1_cm_nx535), .A2 (
          chipmulties_1_cm_nx589), .B0 (B_1__1), .B1 (chipmulties_1_cm_nx573), .B2 (
          chipmulties_1_cm_nx591)) ;
    aoi22 chipmulties_1_cm_ix588 (.Y (chipmulties_1_cm_nx587), .A0 (
          chipmulties_1_cm_nx562), .A1 (chipmulties_1_cm_nx571), .B0 (
          chipmulties_1_cm_nx573), .B1 (chipmulties_1_cm_nx130)) ;
    aoi21 chipmulties_1_cm_ix590 (.Y (chipmulties_1_cm_nx589), .A0 (A_1__2), .A1 (
          A_1__1), .B0 (B_1__4)) ;
    oai21 chipmulties_1_cm_ix592 (.Y (chipmulties_1_cm_nx591), .A0 (
          chipmulties_1_cm_nx46), .A1 (chipmulties_1_cm_nx528), .B0 (A_1__3)) ;
    inv01 chipmulties_1_cm_ix79 (.Y (chipmulties_1_cm_nx78), .A (
          chipmulties_1_cm_nx535)) ;
    inv01 chipmulties_1_cm_ix584 (.Y (chipmulties_1_cm_nx583), .A (
          chipmulties_1_cm_nx46)) ;
    inv01 chipmulties_1_cm_ix23 (.Y (chipmulties_1_cm_nx22), .A (
          chipmulties_1_cm_nx511)) ;
    inv01 chipmulties_1_cm_ix19 (.Y (chipmulties_1_cm_nx18), .A (
          chipmulties_1_cm_nx513)) ;
    inv01 chipmulties_1_cm_ix572 (.Y (chipmulties_1_cm_nx571), .A (
          chipmulties_1_cm_nx2)) ;
    nor02ii chipmulties_1_cm_ix512 (.Y (chipmulties_1_cm_nx511), .A0 (A_1__4), .A1 (
            A_1__3)) ;
    and03 chipmulties_1_cm_ix519 (.Y (chipmulties_1_cm_nx518), .A0 (A_1__3), .A1 (
          chipmulties_1_cm_nx573), .A2 (A_1__1)) ;
    nor02ii chipmulties_1_cm_ix131 (.Y (chipmulties_1_cm_nx130), .A0 (A_1__3), .A1 (
            B_1__1)) ;
    nor04 chipmulties_0_cm_ix41 (.Y (C_0__0), .A0 (chipmulties_0_cm_nx501), .A1 (
          chipmulties_0_cm_nx503), .A2 (chipmulties_0_cm_nx508), .A3 (
          chipmulties_0_cm_nx518)) ;
    inv01 chipmulties_0_cm_ix502 (.Y (chipmulties_0_cm_nx501), .A (A_0__0)) ;
    oai21 chipmulties_0_cm_ix504 (.Y (chipmulties_0_cm_nx503), .A0 (
          chipmulties_0_cm_nx2), .A1 (A_0__2), .B0 (B_0__0)) ;
    nand02 chipmulties_0_cm_ix3 (.Y (chipmulties_0_cm_nx2), .A0 (
           chipmulties_0_cm_nx506), .A1 (A_0__4)) ;
    inv01 chipmulties_0_cm_ix507 (.Y (chipmulties_0_cm_nx506), .A (A_0__3)) ;
    oai21 chipmulties_0_cm_ix509 (.Y (chipmulties_0_cm_nx508), .A0 (
          chipmulties_0_cm_nx2), .A1 (A_0__1), .B0 (chipmulties_0_cm_nx28)) ;
    aoi21 chipmulties_0_cm_ix29 (.Y (chipmulties_0_cm_nx28), .A0 (
          chipmulties_0_cm_nx511), .A1 (A_0__2), .B0 (chipmulties_0_cm_nx513)) ;
    nand03 chipmulties_0_cm_ix514 (.Y (chipmulties_0_cm_nx513), .A0 (
           chipmulties_0_cm_nx10), .A1 (chipmulties_0_cm_nx12), .A2 (
           chipmulties_0_cm_nx14)) ;
    xnor2 chipmulties_0_cm_ix11 (.Y (chipmulties_0_cm_nx10), .A0 (B_0__3), .A1 (
          B_0__4)) ;
    xnor2 chipmulties_0_cm_ix13 (.Y (chipmulties_0_cm_nx12), .A0 (B_0__2), .A1 (
          B_0__1)) ;
    xnor2 chipmulties_0_cm_ix15 (.Y (chipmulties_0_cm_nx14), .A0 (B_0__3), .A1 (
          B_0__2)) ;
    nor02 chipmulties_0_cm_ix75 (.Y (C_0__1), .A0 (chipmulties_0_cm_nx503), .A1 (
          chipmulties_0_cm_nx523)) ;
    aoi32 chipmulties_0_cm_ix524 (.Y (chipmulties_0_cm_nx523), .A0 (
          chipmulties_0_cm_nx52), .A1 (chipmulties_0_cm_nx54), .A2 (
          chipmulties_0_cm_nx28), .B0 (chipmulties_0_cm_nx46), .B1 (
          chipmulties_0_cm_nx68)) ;
    nor02 chipmulties_0_cm_ix53 (.Y (chipmulties_0_cm_nx52), .A0 (B_0__1), .A1 (
          chipmulties_0_cm_nx46)) ;
    nand02 chipmulties_0_cm_ix47 (.Y (chipmulties_0_cm_nx46), .A0 (A_0__0), .A1 (
           A_0__1)) ;
    nand02 chipmulties_0_cm_ix55 (.Y (chipmulties_0_cm_nx54), .A0 (
           chipmulties_0_cm_nx511), .A1 (chipmulties_0_cm_nx528)) ;
    inv01 chipmulties_0_cm_ix529 (.Y (chipmulties_0_cm_nx528), .A (B_0__4)) ;
    ao32 chipmulties_0_cm_ix69 (.Y (chipmulties_0_cm_nx68), .A0 (B_0__1), .A1 (
         A_0__0), .A2 (chipmulties_0_cm_nx62), .B0 (A_0__1), .B1 (
         chipmulties_0_cm_nx28)) ;
    aoi21 chipmulties_0_cm_ix63 (.Y (chipmulties_0_cm_nx62), .A0 (
          chipmulties_0_cm_nx511), .A1 (chipmulties_0_cm_nx528), .B0 (
          chipmulties_0_cm_nx508)) ;
    nor04 chipmulties_0_cm_ix109 (.Y (C_0__2), .A0 (chipmulties_0_cm_nx508), .A1 (
          chipmulties_0_cm_nx533), .A2 (chipmulties_0_cm_nx535), .A3 (
          chipmulties_0_cm_nx537)) ;
    inv01 chipmulties_0_cm_ix534 (.Y (chipmulties_0_cm_nx533), .A (B_0__0)) ;
    nor03 chipmulties_0_cm_ix536 (.Y (chipmulties_0_cm_nx535), .A0 (A_0__0), .A1 (
          A_0__1), .A2 (A_0__2)) ;
    ao22 chipmulties_0_cm_ix538 (.Y (chipmulties_0_cm_nx537), .A0 (
         chipmulties_0_cm_nx539), .A1 (chipmulties_0_cm_nx543), .B0 (
         chipmulties_0_cm_nx545), .B1 (chipmulties_0_cm_nx547)) ;
    oai21 chipmulties_0_cm_ix540 (.Y (chipmulties_0_cm_nx539), .A0 (A_0__2), .A1 (
          B_0__1), .B0 (chipmulties_0_cm_nx541)) ;
    nor02 chipmulties_0_cm_ix542 (.Y (chipmulties_0_cm_nx541), .A0 (A_0__0), .A1 (
          A_0__1)) ;
    xnor2 chipmulties_0_cm_ix544 (.Y (chipmulties_0_cm_nx543), .A0 (B_0__1), .A1 (
          A_0__2)) ;
    oai22 chipmulties_0_cm_ix546 (.Y (chipmulties_0_cm_nx545), .A0 (
          chipmulties_0_cm_nx2), .A1 (chipmulties_0_cm_nx528), .B0 (
          chipmulties_0_cm_nx506), .B1 (A_0__4)) ;
    nand03 chipmulties_0_cm_ix548 (.Y (chipmulties_0_cm_nx547), .A0 (
           chipmulties_0_cm_nx2), .A1 (B_0__4), .A2 (chipmulties_0_cm_nx46)) ;
    aoi21 chipmulties_0_cm_ix185 (.Y (C_0__3), .A0 (chipmulties_0_cm_nx550), .A1 (
          chipmulties_0_cm_nx569), .B0 (chipmulties_0_cm_nx575)) ;
    oai21 chipmulties_0_cm_ix551 (.Y (chipmulties_0_cm_nx550), .A0 (
          chipmulties_0_cm_nx2), .A1 (A_0__1), .B0 (chipmulties_0_cm_nx178)) ;
    oai22 chipmulties_0_cm_ix179 (.Y (chipmulties_0_cm_nx178), .A0 (
          chipmulties_0_cm_nx553), .A1 (chipmulties_0_cm_nx557), .B0 (
          chipmulties_0_cm_nx528), .B1 (chipmulties_0_cm_nx566)) ;
    aoi21 chipmulties_0_cm_ix554 (.Y (chipmulties_0_cm_nx553), .A0 (
          chipmulties_0_cm_nx555), .A1 (chipmulties_0_cm_nx46), .B0 (A_0__4)) ;
    inv01 chipmulties_0_cm_ix556 (.Y (chipmulties_0_cm_nx555), .A (A_0__2)) ;
    nand02 chipmulties_0_cm_ix558 (.Y (chipmulties_0_cm_nx557), .A0 (
           chipmulties_0_cm_nx528), .A1 (chipmulties_0_cm_nx154)) ;
    oai21 chipmulties_0_cm_ix155 (.Y (chipmulties_0_cm_nx154), .A0 (
          chipmulties_0_cm_nx506), .A1 (A_0__0), .B0 (chipmulties_0_cm_nx560)) ;
    aoi22 chipmulties_0_cm_ix561 (.Y (chipmulties_0_cm_nx560), .A0 (
          chipmulties_0_cm_nx562), .A1 (A_0__3), .B0 (chipmulties_0_cm_nx78), .B1 (
          chipmulties_0_cm_nx130)) ;
    inv01 chipmulties_0_cm_ix563 (.Y (chipmulties_0_cm_nx562), .A (B_0__1)) ;
    aoi32 chipmulties_0_cm_ix567 (.Y (chipmulties_0_cm_nx566), .A0 (
          chipmulties_0_cm_nx164), .A1 (chipmulties_0_cm_nx78), .A2 (
          chipmulties_0_cm_nx130), .B0 (A_0__3), .B1 (chipmulties_0_cm_nx541)) ;
    nand02 chipmulties_0_cm_ix165 (.Y (chipmulties_0_cm_nx164), .A0 (
           chipmulties_0_cm_nx555), .A1 (A_0__4)) ;
    or04 chipmulties_0_cm_ix570 (.Y (chipmulties_0_cm_nx569), .A0 (
         chipmulties_0_cm_nx528), .A1 (A_0__1), .A2 (chipmulties_0_cm_nx560), .A3 (
         chipmulties_0_cm_nx571)) ;
    inv01 chipmulties_0_cm_ix574 (.Y (chipmulties_0_cm_nx573), .A (A_0__4)) ;
    nand03 chipmulties_0_cm_ix576 (.Y (chipmulties_0_cm_nx575), .A0 (
           chipmulties_0_cm_nx118), .A1 (B_0__0), .A2 (chipmulties_0_cm_nx18)) ;
    nand03 chipmulties_0_cm_ix119 (.Y (chipmulties_0_cm_nx118), .A0 (B_0__4), .A1 (
           A_0__2), .A2 (A_0__3)) ;
    nor02 chipmulties_0_cm_ix233 (.Y (C_0__4), .A0 (chipmulties_0_cm_nx575), .A1 (
          chipmulties_0_cm_nx580)) ;
    aoi21 chipmulties_0_cm_ix581 (.Y (chipmulties_0_cm_nx580), .A0 (B_0__1), .A1 (
          chipmulties_0_cm_nx192), .B0 (chipmulties_0_cm_nx228)) ;
    aoi21 chipmulties_0_cm_ix193 (.Y (chipmulties_0_cm_nx192), .A0 (
          chipmulties_0_cm_nx583), .A1 (B_0__4), .B0 (chipmulties_0_cm_nx22)) ;
    oai33 chipmulties_0_cm_ix229 (.Y (chipmulties_0_cm_nx228), .A0 (
          chipmulties_0_cm_nx587), .A1 (chipmulties_0_cm_nx535), .A2 (
          chipmulties_0_cm_nx589), .B0 (B_0__1), .B1 (chipmulties_0_cm_nx573), .B2 (
          chipmulties_0_cm_nx591)) ;
    aoi22 chipmulties_0_cm_ix588 (.Y (chipmulties_0_cm_nx587), .A0 (
          chipmulties_0_cm_nx562), .A1 (chipmulties_0_cm_nx571), .B0 (
          chipmulties_0_cm_nx573), .B1 (chipmulties_0_cm_nx130)) ;
    aoi21 chipmulties_0_cm_ix590 (.Y (chipmulties_0_cm_nx589), .A0 (A_0__2), .A1 (
          A_0__1), .B0 (B_0__4)) ;
    oai21 chipmulties_0_cm_ix592 (.Y (chipmulties_0_cm_nx591), .A0 (
          chipmulties_0_cm_nx46), .A1 (chipmulties_0_cm_nx528), .B0 (A_0__3)) ;
    inv01 chipmulties_0_cm_ix79 (.Y (chipmulties_0_cm_nx78), .A (
          chipmulties_0_cm_nx535)) ;
    inv01 chipmulties_0_cm_ix584 (.Y (chipmulties_0_cm_nx583), .A (
          chipmulties_0_cm_nx46)) ;
    inv01 chipmulties_0_cm_ix23 (.Y (chipmulties_0_cm_nx22), .A (
          chipmulties_0_cm_nx511)) ;
    inv01 chipmulties_0_cm_ix19 (.Y (chipmulties_0_cm_nx18), .A (
          chipmulties_0_cm_nx513)) ;
    inv01 chipmulties_0_cm_ix572 (.Y (chipmulties_0_cm_nx571), .A (
          chipmulties_0_cm_nx2)) ;
    nor02ii chipmulties_0_cm_ix512 (.Y (chipmulties_0_cm_nx511), .A0 (A_0__4), .A1 (
            A_0__3)) ;
    and03 chipmulties_0_cm_ix519 (.Y (chipmulties_0_cm_nx518), .A0 (A_0__3), .A1 (
          chipmulties_0_cm_nx573), .A2 (A_0__1)) ;
    nor02ii chipmulties_0_cm_ix131 (.Y (chipmulties_0_cm_nx130), .A0 (A_0__3), .A1 (
            B_0__1)) ;
endmodule

