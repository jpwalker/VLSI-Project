-- types_bdy.vhd
-- Jean P. Walker
-- Body of functions used in 
