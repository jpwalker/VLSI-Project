//
// Verilog description for cell accu, 
// Wed May  8 02:01:03 2019
//
// LeonardoSpectrum Level 3, 2011a.4 
//


module accu ( A_15__4, A_15__3, A_15__2, A_15__1, A_15__0, A_14__4, A_14__3, 
              A_14__2, A_14__1, A_14__0, A_13__4, A_13__3, A_13__2, A_13__1, 
              A_13__0, A_12__4, A_12__3, A_12__2, A_12__1, A_12__0, A_11__4, 
              A_11__3, A_11__2, A_11__1, A_11__0, A_10__4, A_10__3, A_10__2, 
              A_10__1, A_10__0, A_9__4, A_9__3, A_9__2, A_9__1, A_9__0, A_8__4, 
              A_8__3, A_8__2, A_8__1, A_8__0, A_7__4, A_7__3, A_7__2, A_7__1, 
              A_7__0, A_6__4, A_6__3, A_6__2, A_6__1, A_6__0, A_5__4, A_5__3, 
              A_5__2, A_5__1, A_5__0, A_4__4, A_4__3, A_4__2, A_4__1, A_4__0, 
              A_3__4, A_3__3, A_3__2, A_3__1, A_3__0, A_2__4, A_2__3, A_2__2, 
              A_2__1, A_2__0, A_1__4, A_1__3, A_1__2, A_1__1, A_1__0, A_0__4, 
              A_0__3, A_0__2, A_0__1, A_0__0, B ) ;

    input A_15__4 ;
    input A_15__3 ;
    input A_15__2 ;
    input A_15__1 ;
    input A_15__0 ;
    input A_14__4 ;
    input A_14__3 ;
    input A_14__2 ;
    input A_14__1 ;
    input A_14__0 ;
    input A_13__4 ;
    input A_13__3 ;
    input A_13__2 ;
    input A_13__1 ;
    input A_13__0 ;
    input A_12__4 ;
    input A_12__3 ;
    input A_12__2 ;
    input A_12__1 ;
    input A_12__0 ;
    input A_11__4 ;
    input A_11__3 ;
    input A_11__2 ;
    input A_11__1 ;
    input A_11__0 ;
    input A_10__4 ;
    input A_10__3 ;
    input A_10__2 ;
    input A_10__1 ;
    input A_10__0 ;
    input A_9__4 ;
    input A_9__3 ;
    input A_9__2 ;
    input A_9__1 ;
    input A_9__0 ;
    input A_8__4 ;
    input A_8__3 ;
    input A_8__2 ;
    input A_8__1 ;
    input A_8__0 ;
    input A_7__4 ;
    input A_7__3 ;
    input A_7__2 ;
    input A_7__1 ;
    input A_7__0 ;
    input A_6__4 ;
    input A_6__3 ;
    input A_6__2 ;
    input A_6__1 ;
    input A_6__0 ;
    input A_5__4 ;
    input A_5__3 ;
    input A_5__2 ;
    input A_5__1 ;
    input A_5__0 ;
    input A_4__4 ;
    input A_4__3 ;
    input A_4__2 ;
    input A_4__1 ;
    input A_4__0 ;
    input A_3__4 ;
    input A_3__3 ;
    input A_3__2 ;
    input A_3__1 ;
    input A_3__0 ;
    input A_2__4 ;
    input A_2__3 ;
    input A_2__2 ;
    input A_2__1 ;
    input A_2__0 ;
    input A_1__4 ;
    input A_1__3 ;
    input A_1__2 ;
    input A_1__1 ;
    input A_1__0 ;
    input A_0__4 ;
    input A_0__3 ;
    input A_0__2 ;
    input A_0__1 ;
    input A_0__0 ;
    output [8:0]B ;

    wire nx6, nx20, nx34, nx42, nx50, nx54, nx74, nx88, nx98, nx102, nx110, 
         nx114, nx118, nx120, nx138, nx140, nx158, nx160, nx168, nx200, nx204, 
         nx208, nx216, nx224, nx230, nx232, nx234, nx250, nx264, nx274, nx278, 
         nx286, nx290, nx300, nx316, nx330, nx338, nx346, nx350, nx352, nx354, 
         nx372, nx374, nx392, nx394, nx402, nx434, nx438, nx442, nx450, nx458, 
         nx464, nx466, nx468, nx476, nx486, nx488, nx496, nx516, nx518, nx526, 
         nx528, nx548, nx552, nx560, nx568, nx576, nx580, nx582, nx600, nx614, 
         nx624, nx628, nx636, nx640, nx650, nx666, nx680, nx688, nx696, nx700, 
         nx702, nx704, nx722, nx724, nx742, nx744, nx752, nx784, nx788, nx792, 
         nx800, nx808, nx814, nx822, nx824, nx826, nx840, nx854, nx862, nx870, 
         nx874, nx892, nx906, nx916, nx920, nx928, nx932, nx940, nx942, nx944, 
         nx962, nx964, nx972, nx1004, nx1008, nx1012, nx1020, nx1040, nx1042, 
         nx1050, nx1070, nx1072, nx1080, nx1082, nx1102, nx1106, nx1114, nx1122, 
         nx1134, nx1136, nx1138, nx1142, nx1144, nx1156, nx1158, nx1176, nx1178, 
         nx1186, nx1206, nx1208, nx1228, nx1236, nx1240, nx1248, nx1256, nx1272, 
         nx1274, nx1280, nx711, nx713, nx715, nx717, nx719, nx721, nx723, nx725, 
         nx727, nx729, nx731, nx733, nx735, nx737, nx739, nx741, nx743, nx745, 
         nx747, nx749, nx751, nx753, nx759, nx765, nx771, nx773, nx775, nx777, 
         nx779, nx785, nx787, nx789, nx791, nx793, nx799, nx805, nx807, nx809, 
         nx811, nx813, nx819, nx821, nx823, nx825, nx827, nx831, nx833, nx835, 
         nx837, nx839, nx845, nx847, nx849, nx851, nx855, nx857, nx859, nx863, 
         nx869, nx871, nx873, nx875, nx879, nx881, nx883, nx887, nx889, nx891, 
         nx893, nx899, nx901, nx903, nx905, nx909, nx911, nx913, nx917, nx923, 
         nx925, nx927, nx929, nx933, nx935, nx937, nx941, nx947, nx949, nx951, 
         nx955, nx957, nx959, nx963, nx969, nx971, nx977, nx979, nx981, nx983, 
         nx987, nx993, nx995, nx1001, nx1003, nx1005, nx1007, nx1011, nx1013, 
         nx1015, nx1019, nx1025, nx1027, nx1033, nx1035, nx1037, nx1039, nx1043, 
         nx1049, nx1051, nx1057, nx1059, nx1063, nx1067, nx1073, nx1075, nx1077, 
         nx1085, nx1087, nx1089, nx1091, nx1093, nx1095, nx1097, nx1099, nx1101, 
         nx1103, nx1105, nx1113, nx1115, nx1117, nx1119, nx1121, nx1123, nx1125, 
         nx1127, nx1129, nx1135, nx1137, nx1139, nx1147, nx1149, nx1151, nx1153, 
         nx1155, nx1157, nx1159, nx1161, nx1163, nx1165, nx1167, nx1175, nx1177, 
         nx1179, nx1181, nx1183, nx1185, nx1187, nx1189, nx1191, nx1195, nx1201, 
         nx1203, nx1205, nx1209, nx1215, nx1229, nx1239, nx1241, nx1245, nx1251, 
         nx1265, nx1279, nx1285, nx1287, nx1289, nx1291, nx1293, nx1295, nx1297, 
         nx1306, nx1308, nx1311, nx1313, nx1315, nx1317, nx1319, nx1322, nx1324, 
         nx1334, nx1336, nx1338, nx1340, nx1342, nx1344, nx1346, nx1349, nx1351, 
         nx1359, nx1361, nx1363, nx1365, nx1367, nx1375, nx1377, nx1381, nx1383, 
         nx1385, nx1387, nx1390, nx1394, nx1402, nx1408, nx1410, nx1413, nx1417, 
         nx1425, nx1432, nx1435, nx1437, nx1441, nx1445, nx1448, nx1450, nx1456, 
         nx1458, nx1461, nx1465, nx1467, nx1473, nx1475, nx1477, nx1479, nx1482, 
         nx1485, nx1489, nx1492, nx1499, nx1501, nx1503, nx1505, nx1507, nx1509, 
         nx1511, nx1513, nx1515, nx1517, nx1519, nx1521, nx1523, nx1525, nx1527, 
         nx1529, nx1535, nx1537, nx1539, nx1541;



    xor2 ix1303 (.Y (B[0]), .A0 (nx711), .A1 (nx733)) ;
    xnor2 ix712 (.Y (nx711), .A0 (nx713), .A1 (nx723)) ;
    xnor2 ix714 (.Y (nx713), .A0 (nx715), .A1 (nx719)) ;
    oai21 ix716 (.Y (nx715), .A0 (A_0__0), .A1 (A_1__0), .B0 (nx717)) ;
    nand02 ix718 (.Y (nx717), .A0 (A_1__0), .A1 (A_0__0)) ;
    oai21 ix720 (.Y (nx719), .A0 (A_2__0), .A1 (A_3__0), .B0 (nx721)) ;
    nand02 ix722 (.Y (nx721), .A0 (A_3__0), .A1 (A_2__0)) ;
    xnor2 ix724 (.Y (nx723), .A0 (nx725), .A1 (nx729)) ;
    oai21 ix726 (.Y (nx725), .A0 (A_4__0), .A1 (A_5__0), .B0 (nx727)) ;
    nand02 ix728 (.Y (nx727), .A0 (A_5__0), .A1 (A_4__0)) ;
    oai21 ix730 (.Y (nx729), .A0 (A_6__0), .A1 (A_7__0), .B0 (nx731)) ;
    nand02 ix732 (.Y (nx731), .A0 (A_7__0), .A1 (A_6__0)) ;
    xnor2 ix734 (.Y (nx733), .A0 (nx735), .A1 (nx745)) ;
    xnor2 ix736 (.Y (nx735), .A0 (nx737), .A1 (nx741)) ;
    oai21 ix738 (.Y (nx737), .A0 (A_8__0), .A1 (A_9__0), .B0 (nx739)) ;
    nand02 ix740 (.Y (nx739), .A0 (A_9__0), .A1 (A_8__0)) ;
    oai21 ix742 (.Y (nx741), .A0 (A_10__0), .A1 (A_11__0), .B0 (nx743)) ;
    nand02 ix744 (.Y (nx743), .A0 (A_11__0), .A1 (A_10__0)) ;
    xnor2 ix746 (.Y (nx745), .A0 (nx747), .A1 (nx751)) ;
    oai21 ix748 (.Y (nx747), .A0 (A_12__0), .A1 (A_13__0), .B0 (nx749)) ;
    nand02 ix750 (.Y (nx749), .A0 (A_13__0), .A1 (A_12__0)) ;
    oai21 ix752 (.Y (nx751), .A0 (A_14__0), .A1 (A_15__0), .B0 (nx753)) ;
    nand02 ix754 (.Y (nx753), .A0 (A_15__0), .A1 (A_14__0)) ;
    xnor2 ix1297 (.Y (B[1]), .A0 (nx1228), .A1 (nx759)) ;
    nor02 ix1229 (.Y (nx1228), .A0 (nx711), .A1 (nx733)) ;
    xnor2 ix760 (.Y (nx759), .A0 (nx1208), .A1 (nx1206)) ;
    xnor2 ix1209 (.Y (nx1208), .A0 (nx1102), .A1 (nx765)) ;
    nor02 ix1103 (.Y (nx1102), .A0 (nx713), .A1 (nx723)) ;
    xnor2 ix766 (.Y (nx765), .A0 (nx1082), .A1 (nx1080)) ;
    xnor2 ix1083 (.Y (nx1082), .A0 (nx1004), .A1 (nx771)) ;
    nor02 ix1005 (.Y (nx1004), .A0 (nx715), .A1 (nx719)) ;
    xnor2 ix772 (.Y (nx771), .A0 (nx773), .A1 (nx777)) ;
    xnor2 ix774 (.Y (nx773), .A0 (nx717), .A1 (nx775)) ;
    xnor2 ix776 (.Y (nx775), .A0 (A_0__1), .A1 (A_1__1)) ;
    xnor2 ix778 (.Y (nx777), .A0 (nx721), .A1 (nx779)) ;
    xnor2 ix780 (.Y (nx779), .A0 (A_2__1), .A1 (A_3__1)) ;
    xnor2 ix1081 (.Y (nx1080), .A0 (nx784), .A1 (nx785)) ;
    nor02 ix785 (.Y (nx784), .A0 (nx725), .A1 (nx729)) ;
    xnor2 ix786 (.Y (nx785), .A0 (nx787), .A1 (nx791)) ;
    xnor2 ix788 (.Y (nx787), .A0 (nx727), .A1 (nx789)) ;
    xnor2 ix790 (.Y (nx789), .A0 (A_4__1), .A1 (A_5__1)) ;
    xnor2 ix792 (.Y (nx791), .A0 (nx731), .A1 (nx793)) ;
    xnor2 ix794 (.Y (nx793), .A0 (A_6__1), .A1 (A_7__1)) ;
    xnor2 ix1207 (.Y (nx1206), .A0 (nx548), .A1 (nx799)) ;
    nor02 ix549 (.Y (nx548), .A0 (nx735), .A1 (nx745)) ;
    xnor2 ix800 (.Y (nx799), .A0 (nx528), .A1 (nx526)) ;
    xnor2 ix529 (.Y (nx528), .A0 (nx434), .A1 (nx805)) ;
    nor02 ix435 (.Y (nx434), .A0 (nx737), .A1 (nx741)) ;
    xnor2 ix806 (.Y (nx805), .A0 (nx807), .A1 (nx811)) ;
    xnor2 ix808 (.Y (nx807), .A0 (nx739), .A1 (nx809)) ;
    xnor2 ix810 (.Y (nx809), .A0 (A_8__1), .A1 (A_9__1)) ;
    xnor2 ix812 (.Y (nx811), .A0 (nx743), .A1 (nx813)) ;
    xnor2 ix814 (.Y (nx813), .A0 (A_10__1), .A1 (A_11__1)) ;
    xnor2 ix527 (.Y (nx526), .A0 (nx200), .A1 (nx819)) ;
    nor02 ix201 (.Y (nx200), .A0 (nx747), .A1 (nx751)) ;
    xnor2 ix820 (.Y (nx819), .A0 (nx821), .A1 (nx825)) ;
    xnor2 ix822 (.Y (nx821), .A0 (nx749), .A1 (nx823)) ;
    xnor2 ix824 (.Y (nx823), .A0 (A_12__1), .A1 (A_13__1)) ;
    xnor2 ix826 (.Y (nx825), .A0 (nx753), .A1 (nx827)) ;
    xnor2 ix828 (.Y (nx827), .A0 (A_14__1), .A1 (A_15__1)) ;
    xor2 ix1295 (.Y (B[2]), .A0 (nx831), .A1 (nx833)) ;
    mux21 ix832 (.Y (nx831), .A0 (nx1228), .A1 (nx1206), .S0 (nx759)) ;
    xnor2 ix834 (.Y (nx833), .A0 (nx835), .A1 (nx889)) ;
    xnor2 ix836 (.Y (nx835), .A0 (nx837), .A1 (nx839)) ;
    mux21 ix838 (.Y (nx837), .A0 (nx1102), .A1 (nx1080), .S0 (nx765)) ;
    xnor2 ix840 (.Y (nx839), .A0 (nx1072), .A1 (nx1070)) ;
    xnor2 ix1073 (.Y (nx1072), .A0 (nx1008), .A1 (nx847)) ;
    mux21 ix1009 (.Y (nx1008), .A0 (nx845), .A1 (nx777), .S0 (nx771)) ;
    xnor2 ix848 (.Y (nx847), .A0 (nx849), .A1 (nx857)) ;
    xnor2 ix850 (.Y (nx849), .A0 (nx851), .A1 (nx855)) ;
    aoi32 ix852 (.Y (nx851), .A0 (A_1__0), .A1 (A_0__0), .A2 (nx892), .B0 (
          A_0__1), .B1 (A_1__1)) ;
    xnor2 ix856 (.Y (nx855), .A0 (A_0__2), .A1 (A_1__2)) ;
    xnor2 ix858 (.Y (nx857), .A0 (nx859), .A1 (nx863)) ;
    aoi32 ix860 (.Y (nx859), .A0 (A_3__0), .A1 (A_2__0), .A2 (nx840), .B0 (
          A_2__1), .B1 (A_3__1)) ;
    xnor2 ix864 (.Y (nx863), .A0 (A_2__2), .A1 (A_3__2)) ;
    xnor2 ix1071 (.Y (nx1070), .A0 (nx788), .A1 (nx871)) ;
    mux21 ix789 (.Y (nx788), .A0 (nx869), .A1 (nx791), .S0 (nx785)) ;
    xnor2 ix872 (.Y (nx871), .A0 (nx873), .A1 (nx881)) ;
    xnor2 ix874 (.Y (nx873), .A0 (nx875), .A1 (nx879)) ;
    aoi32 ix876 (.Y (nx875), .A0 (A_5__0), .A1 (A_4__0), .A2 (nx666), .B0 (
          A_4__1), .B1 (A_5__1)) ;
    xnor2 ix880 (.Y (nx879), .A0 (A_4__2), .A1 (A_5__2)) ;
    xnor2 ix882 (.Y (nx881), .A0 (nx883), .A1 (nx887)) ;
    aoi32 ix884 (.Y (nx883), .A0 (A_7__0), .A1 (A_6__0), .A2 (nx600), .B0 (
          A_6__1), .B1 (A_7__1)) ;
    xnor2 ix888 (.Y (nx887), .A0 (A_6__2), .A1 (A_7__2)) ;
    xnor2 ix890 (.Y (nx889), .A0 (nx891), .A1 (nx893)) ;
    mux21 ix892 (.Y (nx891), .A0 (nx548), .A1 (nx526), .S0 (nx799)) ;
    xnor2 ix894 (.Y (nx893), .A0 (nx518), .A1 (nx516)) ;
    xnor2 ix519 (.Y (nx518), .A0 (nx438), .A1 (nx901)) ;
    mux21 ix439 (.Y (nx438), .A0 (nx899), .A1 (nx811), .S0 (nx805)) ;
    xnor2 ix902 (.Y (nx901), .A0 (nx903), .A1 (nx911)) ;
    xnor2 ix904 (.Y (nx903), .A0 (nx905), .A1 (nx909)) ;
    aoi32 ix906 (.Y (nx905), .A0 (A_9__0), .A1 (A_8__0), .A2 (nx316), .B0 (
          A_8__1), .B1 (A_9__1)) ;
    xnor2 ix910 (.Y (nx909), .A0 (A_8__2), .A1 (A_9__2)) ;
    xnor2 ix912 (.Y (nx911), .A0 (nx913), .A1 (nx917)) ;
    aoi32 ix914 (.Y (nx913), .A0 (A_11__0), .A1 (A_10__0), .A2 (nx250), .B0 (
          A_10__1), .B1 (A_11__1)) ;
    xnor2 ix918 (.Y (nx917), .A0 (A_10__2), .A1 (A_11__2)) ;
    xnor2 ix517 (.Y (nx516), .A0 (nx204), .A1 (nx925)) ;
    mux21 ix205 (.Y (nx204), .A0 (nx923), .A1 (nx825), .S0 (nx819)) ;
    xnor2 ix926 (.Y (nx925), .A0 (nx927), .A1 (nx935)) ;
    xnor2 ix928 (.Y (nx927), .A0 (nx929), .A1 (nx933)) ;
    aoi32 ix930 (.Y (nx929), .A0 (A_13__0), .A1 (A_12__0), .A2 (nx74), .B0 (
          A_12__1), .B1 (A_13__1)) ;
    xnor2 ix934 (.Y (nx933), .A0 (A_12__2), .A1 (A_13__2)) ;
    xnor2 ix936 (.Y (nx935), .A0 (nx937), .A1 (nx941)) ;
    aoi32 ix938 (.Y (nx937), .A0 (A_15__0), .A1 (A_14__0), .A2 (nx20), .B0 (
          A_14__1), .B1 (A_15__1)) ;
    xnor2 ix942 (.Y (nx941), .A0 (A_14__2), .A1 (A_15__2)) ;
    xnor2 ix1293 (.Y (B[3]), .A0 (nx1236), .A1 (nx947)) ;
    mux21 ix1237 (.Y (nx1236), .A0 (nx831), .A1 (nx889), .S0 (nx833)) ;
    xnor2 ix948 (.Y (nx947), .A0 (nx949), .A1 (nx1005)) ;
    xnor2 ix950 (.Y (nx949), .A0 (nx951), .A1 (nx955)) ;
    mux21 ix952 (.Y (nx951), .A0 (nx1106), .A1 (nx1070), .S0 (nx839)) ;
    xnor2 ix956 (.Y (nx955), .A0 (nx957), .A1 (nx981)) ;
    xnor2 ix958 (.Y (nx957), .A0 (nx959), .A1 (nx963)) ;
    mux21 ix960 (.Y (nx959), .A0 (nx1008), .A1 (nx972), .S0 (nx847)) ;
    xnor2 ix964 (.Y (nx963), .A0 (nx964), .A1 (nx962)) ;
    xnor2 ix965 (.Y (nx964), .A0 (nx906), .A1 (nx971)) ;
    mux21 ix907 (.Y (nx906), .A0 (nx851), .A1 (nx969), .S0 (nx855)) ;
    inv01 ix970 (.Y (nx969), .A (A_0__2)) ;
    xnor2 ix972 (.Y (nx971), .A0 (A_0__3), .A1 (A_1__3)) ;
    xnor2 ix963 (.Y (nx962), .A0 (nx854), .A1 (nx979)) ;
    mux21 ix855 (.Y (nx854), .A0 (nx859), .A1 (nx977), .S0 (nx863)) ;
    inv01 ix978 (.Y (nx977), .A (A_2__2)) ;
    xnor2 ix980 (.Y (nx979), .A0 (A_2__3), .A1 (A_3__3)) ;
    xnor2 ix982 (.Y (nx981), .A0 (nx983), .A1 (nx987)) ;
    mux21 ix984 (.Y (nx983), .A0 (nx788), .A1 (nx752), .S0 (nx871)) ;
    xnor2 ix988 (.Y (nx987), .A0 (nx744), .A1 (nx742)) ;
    xnor2 ix745 (.Y (nx744), .A0 (nx680), .A1 (nx995)) ;
    mux21 ix681 (.Y (nx680), .A0 (nx875), .A1 (nx993), .S0 (nx879)) ;
    inv01 ix994 (.Y (nx993), .A (A_4__2)) ;
    xnor2 ix996 (.Y (nx995), .A0 (A_4__3), .A1 (A_5__3)) ;
    xnor2 ix743 (.Y (nx742), .A0 (nx614), .A1 (nx1003)) ;
    mux21 ix615 (.Y (nx614), .A0 (nx883), .A1 (nx1001), .S0 (nx887)) ;
    inv01 ix1002 (.Y (nx1001), .A (A_6__2)) ;
    xnor2 ix1004 (.Y (nx1003), .A0 (A_6__3), .A1 (A_7__3)) ;
    xnor2 ix1006 (.Y (nx1005), .A0 (nx1007), .A1 (nx1011)) ;
    mux21 ix1008 (.Y (nx1007), .A0 (nx552), .A1 (nx516), .S0 (nx893)) ;
    xnor2 ix1012 (.Y (nx1011), .A0 (nx1013), .A1 (nx1037)) ;
    xnor2 ix1014 (.Y (nx1013), .A0 (nx1015), .A1 (nx1019)) ;
    mux21 ix1016 (.Y (nx1015), .A0 (nx438), .A1 (nx402), .S0 (nx901)) ;
    xnor2 ix1020 (.Y (nx1019), .A0 (nx394), .A1 (nx392)) ;
    xnor2 ix395 (.Y (nx394), .A0 (nx330), .A1 (nx1027)) ;
    mux21 ix331 (.Y (nx330), .A0 (nx905), .A1 (nx1025), .S0 (nx909)) ;
    inv01 ix1026 (.Y (nx1025), .A (A_8__2)) ;
    xnor2 ix1028 (.Y (nx1027), .A0 (A_8__3), .A1 (A_9__3)) ;
    xnor2 ix393 (.Y (nx392), .A0 (nx264), .A1 (nx1035)) ;
    mux21 ix265 (.Y (nx264), .A0 (nx913), .A1 (nx1033), .S0 (nx917)) ;
    inv01 ix1034 (.Y (nx1033), .A (A_10__2)) ;
    xnor2 ix1036 (.Y (nx1035), .A0 (A_10__3), .A1 (A_11__3)) ;
    xnor2 ix1038 (.Y (nx1037), .A0 (nx1039), .A1 (nx1043)) ;
    mux21 ix1040 (.Y (nx1039), .A0 (nx204), .A1 (nx168), .S0 (nx925)) ;
    xnor2 ix1044 (.Y (nx1043), .A0 (nx160), .A1 (nx158)) ;
    xnor2 ix161 (.Y (nx160), .A0 (nx88), .A1 (nx1051)) ;
    mux21 ix89 (.Y (nx88), .A0 (nx929), .A1 (nx1049), .S0 (nx933)) ;
    inv01 ix1050 (.Y (nx1049), .A (A_12__2)) ;
    xnor2 ix1052 (.Y (nx1051), .A0 (A_12__3), .A1 (A_13__3)) ;
    xnor2 ix159 (.Y (nx158), .A0 (nx34), .A1 (nx1059)) ;
    mux21 ix35 (.Y (nx34), .A0 (nx937), .A1 (nx1057), .S0 (nx941)) ;
    inv01 ix1058 (.Y (nx1057), .A (A_14__2)) ;
    xnor2 ix1060 (.Y (nx1059), .A0 (A_14__3), .A1 (A_15__3)) ;
    xor2 ix1291 (.Y (B[4]), .A0 (nx1063), .A1 (nx1067)) ;
    mux21 ix1064 (.Y (nx1063), .A0 (nx1236), .A1 (nx1186), .S0 (nx947)) ;
    xnor2 ix1068 (.Y (nx1067), .A0 (nx1178), .A1 (nx1176)) ;
    xnor2 ix1179 (.Y (nx1178), .A0 (nx1114), .A1 (nx1073)) ;
    mux21 ix1115 (.Y (nx1114), .A0 (nx951), .A1 (nx981), .S0 (nx955)) ;
    xnor2 ix1074 (.Y (nx1073), .A0 (nx1075), .A1 (nx1103)) ;
    xnor2 ix1076 (.Y (nx1075), .A0 (nx1077), .A1 (nx1085)) ;
    mux21 ix1078 (.Y (nx1077), .A0 (nx1012), .A1 (nx962), .S0 (nx963)) ;
    xnor2 ix1086 (.Y (nx1085), .A0 (nx1087), .A1 (nx1095)) ;
    mux21 ix1090 (.Y (nx1089), .A0 (nx906), .A1 (A_0__3), .S0 (nx971)) ;
    oai21 ix1092 (.Y (nx1091), .A0 (A_0__4), .A1 (A_1__4), .B0 (nx1093)) ;
    nand02 ix1094 (.Y (nx1093), .A0 (A_1__4), .A1 (A_0__4)) ;
    mux21 ix1098 (.Y (nx1097), .A0 (nx854), .A1 (A_2__3), .S0 (nx979)) ;
    oai21 ix1100 (.Y (nx1099), .A0 (A_2__4), .A1 (A_3__4), .B0 (nx1101)) ;
    nand02 ix1102 (.Y (nx1101), .A0 (A_3__4), .A1 (A_2__4)) ;
    xnor2 ix1104 (.Y (nx1103), .A0 (nx1105), .A1 (nx1113)) ;
    mux21 ix1106 (.Y (nx1105), .A0 (nx792), .A1 (nx742), .S0 (nx987)) ;
    xnor2 ix1114 (.Y (nx1113), .A0 (nx1115), .A1 (nx1123)) ;
    mux21 ix1118 (.Y (nx1117), .A0 (nx680), .A1 (A_4__3), .S0 (nx995)) ;
    oai21 ix1120 (.Y (nx1119), .A0 (A_4__4), .A1 (A_5__4), .B0 (nx1121)) ;
    nand02 ix1122 (.Y (nx1121), .A0 (A_5__4), .A1 (A_4__4)) ;
    mux21 ix1126 (.Y (nx1125), .A0 (nx614), .A1 (A_6__3), .S0 (nx1003)) ;
    oai21 ix1128 (.Y (nx1127), .A0 (A_6__4), .A1 (A_7__4), .B0 (nx1129)) ;
    nand02 ix1130 (.Y (nx1129), .A0 (A_7__4), .A1 (A_6__4)) ;
    xnor2 ix1177 (.Y (nx1176), .A0 (nx560), .A1 (nx1135)) ;
    mux21 ix561 (.Y (nx560), .A0 (nx1007), .A1 (nx1037), .S0 (nx1011)) ;
    xnor2 ix1136 (.Y (nx1135), .A0 (nx1137), .A1 (nx1165)) ;
    xnor2 ix1138 (.Y (nx1137), .A0 (nx1139), .A1 (nx1147)) ;
    mux21 ix1140 (.Y (nx1139), .A0 (nx442), .A1 (nx392), .S0 (nx1019)) ;
    xnor2 ix1148 (.Y (nx1147), .A0 (nx1149), .A1 (nx1157)) ;
    mux21 ix1152 (.Y (nx1151), .A0 (nx330), .A1 (A_8__3), .S0 (nx1027)) ;
    oai21 ix1154 (.Y (nx1153), .A0 (A_8__4), .A1 (A_9__4), .B0 (nx1155)) ;
    nand02 ix1156 (.Y (nx1155), .A0 (A_9__4), .A1 (A_8__4)) ;
    mux21 ix1160 (.Y (nx1159), .A0 (nx264), .A1 (A_10__3), .S0 (nx1035)) ;
    oai21 ix1162 (.Y (nx1161), .A0 (A_10__4), .A1 (A_11__4), .B0 (nx1163)) ;
    nand02 ix1164 (.Y (nx1163), .A0 (A_11__4), .A1 (A_10__4)) ;
    xnor2 ix1166 (.Y (nx1165), .A0 (nx1167), .A1 (nx1175)) ;
    mux21 ix1168 (.Y (nx1167), .A0 (nx208), .A1 (nx158), .S0 (nx1043)) ;
    xnor2 ix1176 (.Y (nx1175), .A0 (nx1177), .A1 (nx1185)) ;
    mux21 ix1180 (.Y (nx1179), .A0 (nx88), .A1 (A_12__3), .S0 (nx1051)) ;
    oai21 ix1182 (.Y (nx1181), .A0 (A_12__4), .A1 (A_13__4), .B0 (nx1183)) ;
    nand02 ix1184 (.Y (nx1183), .A0 (A_13__4), .A1 (A_12__4)) ;
    mux21 ix1188 (.Y (nx1187), .A0 (nx34), .A1 (A_14__3), .S0 (nx1059)) ;
    oai21 ix1190 (.Y (nx1189), .A0 (A_14__4), .A1 (A_15__4), .B0 (nx1191)) ;
    nand02 ix1192 (.Y (nx1191), .A0 (A_15__4), .A1 (A_14__4)) ;
    xor2 ix1289 (.Y (B[5]), .A0 (nx1195), .A1 (nx1201)) ;
    mux21 ix1196 (.Y (nx1195), .A0 (nx1240), .A1 (nx1176), .S0 (nx1067)) ;
    xnor2 ix1202 (.Y (nx1201), .A0 (nx1203), .A1 (nx1239)) ;
    xnor2 ix1204 (.Y (nx1203), .A0 (nx1205), .A1 (nx1209)) ;
    mux21 ix1206 (.Y (nx1205), .A0 (nx1114), .A1 (nx1050), .S0 (nx1073)) ;
    xnor2 ix1210 (.Y (nx1209), .A0 (nx1042), .A1 (nx1040)) ;
    xnor2 ix1043 (.Y (nx1042), .A0 (nx1020), .A1 (nx1215)) ;
    mux21 ix1021 (.Y (nx1020), .A0 (nx1077), .A1 (nx1095), .S0 (nx1085)) ;
    xnor2 ix1216 (.Y (nx1215), .A0 (nx944), .A1 (nx942)) ;
    oai21 ix921 (.Y (nx920), .A0 (nx1089), .A1 (nx1499), .B0 (nx1093)) ;
    oai21 ix863 (.Y (nx862), .A0 (nx1503), .A1 (nx1097), .B0 (nx1101)) ;
    xnor2 ix1041 (.Y (nx1040), .A0 (nx800), .A1 (nx1229)) ;
    mux21 ix801 (.Y (nx800), .A0 (nx1105), .A1 (nx1123), .S0 (nx1113)) ;
    xnor2 ix1230 (.Y (nx1229), .A0 (nx724), .A1 (nx722)) ;
    oai21 ix689 (.Y (nx688), .A0 (nx1507), .A1 (nx1117), .B0 (nx1121)) ;
    oai21 ix629 (.Y (nx628), .A0 (nx1125), .A1 (nx1511), .B0 (nx1129)) ;
    xnor2 ix1240 (.Y (nx1239), .A0 (nx1241), .A1 (nx1245)) ;
    mux21 ix1242 (.Y (nx1241), .A0 (nx560), .A1 (nx496), .S0 (nx1135)) ;
    xnor2 ix1246 (.Y (nx1245), .A0 (nx488), .A1 (nx486)) ;
    xnor2 ix489 (.Y (nx488), .A0 (nx450), .A1 (nx1251)) ;
    mux21 ix451 (.Y (nx450), .A0 (nx1139), .A1 (nx1157), .S0 (nx1147)) ;
    xnor2 ix1252 (.Y (nx1251), .A0 (nx374), .A1 (nx372)) ;
    oai21 ix339 (.Y (nx338), .A0 (nx1515), .A1 (nx1151), .B0 (nx1155)) ;
    oai21 ix279 (.Y (nx278), .A0 (nx1159), .A1 (nx1519), .B0 (nx1163)) ;
    xnor2 ix487 (.Y (nx486), .A0 (nx216), .A1 (nx1265)) ;
    mux21 ix217 (.Y (nx216), .A0 (nx1167), .A1 (nx1185), .S0 (nx1175)) ;
    xnor2 ix1266 (.Y (nx1265), .A0 (nx140), .A1 (nx138)) ;
    oai21 ix103 (.Y (nx102), .A0 (nx1179), .A1 (nx1523), .B0 (nx1183)) ;
    oai21 ix43 (.Y (nx42), .A0 (nx1527), .A1 (nx1187), .B0 (nx1191)) ;
    xnor2 ix1287 (.Y (B[6]), .A0 (nx1248), .A1 (nx1279)) ;
    mux21 ix1249 (.Y (nx1248), .A0 (nx1195), .A1 (nx1239), .S0 (nx1201)) ;
    xnor2 ix1280 (.Y (nx1279), .A0 (nx1158), .A1 (nx1156)) ;
    xnor2 ix1159 (.Y (nx1158), .A0 (nx1122), .A1 (nx1287)) ;
    mux21 ix1123 (.Y (nx1122), .A0 (nx1205), .A1 (nx1285), .S0 (nx1209)) ;
    xnor2 ix1288 (.Y (nx1287), .A0 (nx1289), .A1 (nx1311)) ;
    xnor2 ix1290 (.Y (nx1289), .A0 (nx1291), .A1 (nx1293)) ;
    mux21 ix1292 (.Y (nx1291), .A0 (nx1020), .A1 (nx942), .S0 (nx1215)) ;
    xnor2 ix1294 (.Y (nx1293), .A0 (nx1295), .A1 (nx1306)) ;
    aoi22 ix1298 (.Y (nx1297), .A0 (A_1__4), .A1 (A_0__4), .B0 (nx920), .B1 (
          nx916)) ;
    aoi22 ix1309 (.Y (nx1308), .A0 (A_3__4), .A1 (A_2__4), .B0 (nx1541), .B1 (
          nx862)) ;
    xnor2 ix1312 (.Y (nx1311), .A0 (nx1313), .A1 (nx1315)) ;
    mux21 ix1314 (.Y (nx1313), .A0 (nx800), .A1 (nx722), .S0 (nx1229)) ;
    xnor2 ix1316 (.Y (nx1315), .A0 (nx1317), .A1 (nx1322)) ;
    aoi22 ix1320 (.Y (nx1319), .A0 (A_5__4), .A1 (A_4__4), .B0 (nx1539), .B1 (
          nx688)) ;
    aoi22 ix1325 (.Y (nx1324), .A0 (A_7__4), .A1 (A_6__4), .B0 (nx628), .B1 (
          nx624)) ;
    xnor2 ix1157 (.Y (nx1156), .A0 (nx568), .A1 (nx1336)) ;
    mux21 ix569 (.Y (nx568), .A0 (nx1241), .A1 (nx1334), .S0 (nx1245)) ;
    xnor2 ix1337 (.Y (nx1336), .A0 (nx1338), .A1 (nx1359)) ;
    xnor2 ix1339 (.Y (nx1338), .A0 (nx1340), .A1 (nx1342)) ;
    mux21 ix1341 (.Y (nx1340), .A0 (nx450), .A1 (nx372), .S0 (nx1251)) ;
    xnor2 ix1343 (.Y (nx1342), .A0 (nx1344), .A1 (nx1349)) ;
    aoi22 ix1347 (.Y (nx1346), .A0 (A_9__4), .A1 (A_8__4), .B0 (nx1537), .B1 (
          nx338)) ;
    aoi22 ix1352 (.Y (nx1351), .A0 (A_11__4), .A1 (A_10__4), .B0 (nx278), .B1 (
          nx274)) ;
    xnor2 ix1360 (.Y (nx1359), .A0 (nx1361), .A1 (nx1363)) ;
    mux21 ix1362 (.Y (nx1361), .A0 (nx216), .A1 (nx138), .S0 (nx1265)) ;
    xnor2 ix1364 (.Y (nx1363), .A0 (nx1365), .A1 (nx1375)) ;
    aoi22 ix1368 (.Y (nx1367), .A0 (A_13__4), .A1 (A_12__4), .B0 (nx102), .B1 (
          nx98)) ;
    aoi22 ix1378 (.Y (nx1377), .A0 (A_15__4), .A1 (A_14__4), .B0 (nx1535), .B1 (
          nx42)) ;
    xor2 ix1285 (.Y (B[7]), .A0 (nx1381), .A1 (nx1383)) ;
    mux21 ix1382 (.Y (nx1381), .A0 (nx1248), .A1 (nx1156), .S0 (nx1279)) ;
    xnor2 ix1384 (.Y (nx1383), .A0 (nx1385), .A1 (nx1408)) ;
    xnor2 ix1386 (.Y (nx1385), .A0 (nx1387), .A1 (nx1390)) ;
    mux21 ix1388 (.Y (nx1387), .A0 (nx1122), .A1 (nx940), .S0 (nx1287)) ;
    xnor2 ix1391 (.Y (nx1390), .A0 (nx1142), .A1 (nx1144)) ;
    xnor2 ix1143 (.Y (nx1142), .A0 (nx1134), .A1 (nx1394)) ;
    mux21 ix1135 (.Y (nx1134), .A0 (nx1291), .A1 (nx1306), .S0 (nx1293)) ;
    xnor2 ix1395 (.Y (nx1394), .A0 (nx1136), .A1 (nx1138)) ;
    oai21 ix929 (.Y (nx928), .A0 (nx1297), .A1 (nx1499), .B0 (nx1093)) ;
    oai21 ix871 (.Y (nx870), .A0 (nx1503), .A1 (nx1308), .B0 (nx1101)) ;
    xnor2 ix1145 (.Y (nx1144), .A0 (nx808), .A1 (nx1402)) ;
    mux21 ix809 (.Y (nx808), .A0 (nx1313), .A1 (nx1322), .S0 (nx1315)) ;
    xnor2 ix1403 (.Y (nx1402), .A0 (nx704), .A1 (nx702)) ;
    oai21 ix697 (.Y (nx696), .A0 (nx1507), .A1 (nx1319), .B0 (nx1121)) ;
    oai21 ix637 (.Y (nx636), .A0 (nx1324), .A1 (nx1511), .B0 (nx1129)) ;
    xnor2 ix1409 (.Y (nx1408), .A0 (nx1410), .A1 (nx1413)) ;
    mux21 ix1411 (.Y (nx1410), .A0 (nx568), .A1 (nx476), .S0 (nx1336)) ;
    xnor2 ix1414 (.Y (nx1413), .A0 (nx468), .A1 (nx466)) ;
    xnor2 ix469 (.Y (nx468), .A0 (nx458), .A1 (nx1417)) ;
    mux21 ix459 (.Y (nx458), .A0 (nx1340), .A1 (nx1349), .S0 (nx1342)) ;
    xnor2 ix1418 (.Y (nx1417), .A0 (nx354), .A1 (nx352)) ;
    oai21 ix347 (.Y (nx346), .A0 (nx1515), .A1 (nx1346), .B0 (nx1155)) ;
    oai21 ix287 (.Y (nx286), .A0 (nx1351), .A1 (nx1519), .B0 (nx1163)) ;
    xnor2 ix467 (.Y (nx466), .A0 (nx224), .A1 (nx1425)) ;
    mux21 ix225 (.Y (nx224), .A0 (nx1361), .A1 (nx1375), .S0 (nx1363)) ;
    xnor2 ix1426 (.Y (nx1425), .A0 (nx120), .A1 (nx118)) ;
    oai21 ix111 (.Y (nx110), .A0 (nx1367), .A1 (nx1523), .B0 (nx1183)) ;
    oai21 ix51 (.Y (nx50), .A0 (nx1527), .A1 (nx1377), .B0 (nx1191)) ;
    xnor2 ix1283 (.Y (B[8]), .A0 (nx1432), .A1 (nx1280)) ;
    xnor2 ix1433 (.Y (nx1432), .A0 (nx234), .A1 (nx582)) ;
    xnor2 ix235 (.Y (nx234), .A0 (nx1435), .A1 (nx232)) ;
    xnor2 ix1438 (.Y (nx1437), .A0 (nx54), .A1 (A_12__4)) ;
    oai21 ix55 (.Y (nx54), .A0 (nx1529), .A1 (nx1377), .B0 (nx1191)) ;
    xnor2 ix233 (.Y (nx232), .A0 (nx1441), .A1 (nx230)) ;
    xnor2 ix1442 (.Y (nx1441), .A0 (A_13__4), .A1 (nx114)) ;
    oai21 ix115 (.Y (nx114), .A0 (nx1367), .A1 (nx1525), .B0 (nx1183)) ;
    xnor2 ix231 (.Y (nx230), .A0 (nx1445), .A1 (A_10__4)) ;
    mux21 ix1446 (.Y (nx1445), .A0 (nx224), .A1 (nx118), .S0 (nx1425)) ;
    xnor2 ix583 (.Y (nx582), .A0 (nx1448), .A1 (nx580)) ;
    xnor2 ix1451 (.Y (nx1450), .A0 (A_11__4), .A1 (nx290)) ;
    oai21 ix291 (.Y (nx290), .A0 (nx1351), .A1 (nx1521), .B0 (nx1163)) ;
    xnor2 ix581 (.Y (nx580), .A0 (nx464), .A1 (nx1458)) ;
    xnor2 ix465 (.Y (nx464), .A0 (nx350), .A1 (nx1456)) ;
    oai21 ix351 (.Y (nx350), .A0 (nx1517), .A1 (nx1346), .B0 (nx1155)) ;
    mux21 ix1457 (.Y (nx1456), .A0 (nx458), .A1 (nx352), .S0 (nx1417)) ;
    xnor2 ix1459 (.Y (nx1458), .A0 (nx576), .A1 (A_6__4)) ;
    mux21 ix577 (.Y (nx576), .A0 (nx1410), .A1 (nx1461), .S0 (nx1413)) ;
    xnor2 ix1281 (.Y (nx1280), .A0 (nx826), .A1 (nx1475)) ;
    xnor2 ix827 (.Y (nx826), .A0 (nx1465), .A1 (nx824)) ;
    xnor2 ix1468 (.Y (nx1467), .A0 (A_7__4), .A1 (nx640)) ;
    oai21 ix641 (.Y (nx640), .A0 (nx1324), .A1 (nx1513), .B0 (nx1129)) ;
    xnor2 ix815 (.Y (nx814), .A0 (nx700), .A1 (nx1473)) ;
    oai21 ix701 (.Y (nx700), .A0 (nx1509), .A1 (nx1319), .B0 (nx1121)) ;
    mux21 ix1474 (.Y (nx1473), .A0 (nx808), .A1 (nx702), .S0 (nx1402)) ;
    xnor2 ix1476 (.Y (nx1475), .A0 (nx1477), .A1 (nx1485)) ;
    xnor2 ix1478 (.Y (nx1477), .A0 (nx1479), .A1 (nx1482)) ;
    xnor2 ix1480 (.Y (nx1479), .A0 (nx874), .A1 (A_0__4)) ;
    oai21 ix875 (.Y (nx874), .A0 (nx1505), .A1 (nx1308), .B0 (nx1101)) ;
    xnor2 ix1483 (.Y (nx1482), .A0 (A_1__4), .A1 (nx932)) ;
    oai21 ix933 (.Y (nx932), .A0 (nx1297), .A1 (nx1501), .B0 (nx1093)) ;
    xnor2 ix1486 (.Y (nx1485), .A0 (nx1256), .A1 (nx1274)) ;
    mux21 ix1257 (.Y (nx1256), .A0 (nx1381), .A1 (nx1408), .S0 (nx1383)) ;
    xnor2 ix1275 (.Y (nx1274), .A0 (nx1489), .A1 (nx1272)) ;
    mux21 ix1490 (.Y (nx1489), .A0 (nx1134), .A1 (nx1138), .S0 (nx1394)) ;
    mux21 ix1273 (.Y (nx1272), .A0 (nx1387), .A1 (nx1492), .S0 (nx1390)) ;
    inv01 ix1241 (.Y (nx1240), .A (nx1063)) ;
    inv01 ix1187 (.Y (nx1186), .A (nx1005)) ;
    inv01 ix1493 (.Y (nx1492), .A (nx1144)) ;
    inv01 ix1107 (.Y (nx1106), .A (nx837)) ;
    inv01 ix1051 (.Y (nx1050), .A (nx1103)) ;
    inv01 ix1286 (.Y (nx1285), .A (nx1040)) ;
    inv01 ix1013 (.Y (nx1012), .A (nx959)) ;
    inv01 ix846 (.Y (nx845), .A (nx1004)) ;
    inv01 ix973 (.Y (nx972), .A (nx857)) ;
    inv01 ix941 (.Y (nx940), .A (nx1311)) ;
    inv01 ix917 (.Y (nx916), .A (nx1091)) ;
    inv01 ix893 (.Y (nx892), .A (nx775)) ;
    inv01 ix841 (.Y (nx840), .A (nx779)) ;
    inv01 ix823 (.Y (nx822), .A (nx1099)) ;
    inv01 ix793 (.Y (nx792), .A (nx983)) ;
    inv01 ix870 (.Y (nx869), .A (nx784)) ;
    inv01 ix753 (.Y (nx752), .A (nx881)) ;
    inv01 ix667 (.Y (nx666), .A (nx789)) ;
    inv01 ix651 (.Y (nx650), .A (nx1119)) ;
    inv01 ix625 (.Y (nx624), .A (nx1127)) ;
    inv01 ix601 (.Y (nx600), .A (nx793)) ;
    inv01 ix553 (.Y (nx552), .A (nx891)) ;
    inv01 ix497 (.Y (nx496), .A (nx1165)) ;
    inv01 ix1335 (.Y (nx1334), .A (nx486)) ;
    inv01 ix477 (.Y (nx476), .A (nx1359)) ;
    inv01 ix1462 (.Y (nx1461), .A (nx466)) ;
    inv01 ix443 (.Y (nx442), .A (nx1015)) ;
    inv01 ix900 (.Y (nx899), .A (nx434)) ;
    inv01 ix403 (.Y (nx402), .A (nx911)) ;
    inv01 ix317 (.Y (nx316), .A (nx809)) ;
    inv01 ix301 (.Y (nx300), .A (nx1153)) ;
    inv01 ix275 (.Y (nx274), .A (nx1161)) ;
    inv01 ix251 (.Y (nx250), .A (nx813)) ;
    inv01 ix209 (.Y (nx208), .A (nx1039)) ;
    inv01 ix924 (.Y (nx923), .A (nx200)) ;
    inv01 ix169 (.Y (nx168), .A (nx935)) ;
    inv01 ix99 (.Y (nx98), .A (nx1181)) ;
    inv01 ix75 (.Y (nx74), .A (nx823)) ;
    inv01 ix21 (.Y (nx20), .A (nx827)) ;
    inv01 ix7 (.Y (nx6), .A (nx1189)) ;
    inv01 ix1498 (.Y (nx1499), .A (nx916)) ;
    inv01 ix1500 (.Y (nx1501), .A (nx916)) ;
    inv01 ix1502 (.Y (nx1503), .A (nx1541)) ;
    inv01 ix1504 (.Y (nx1505), .A (nx1541)) ;
    inv01 ix1506 (.Y (nx1507), .A (nx1539)) ;
    inv01 ix1508 (.Y (nx1509), .A (nx1539)) ;
    inv01 ix1510 (.Y (nx1511), .A (nx624)) ;
    inv01 ix1512 (.Y (nx1513), .A (nx624)) ;
    inv01 ix1514 (.Y (nx1515), .A (nx1537)) ;
    inv01 ix1516 (.Y (nx1517), .A (nx1537)) ;
    inv01 ix1518 (.Y (nx1519), .A (nx274)) ;
    inv01 ix1520 (.Y (nx1521), .A (nx274)) ;
    inv01 ix1522 (.Y (nx1523), .A (nx98)) ;
    inv01 ix1524 (.Y (nx1525), .A (nx98)) ;
    inv01 ix1526 (.Y (nx1527), .A (nx1535)) ;
    inv01 ix1528 (.Y (nx1529), .A (nx1535)) ;
    xor2 ix1088 (.Y (nx1087), .A0 (nx1089), .A1 (nx916)) ;
    xor2 ix1096 (.Y (nx1095), .A0 (nx1097), .A1 (nx1541)) ;
    xor2 ix1116 (.Y (nx1115), .A0 (nx1117), .A1 (nx1539)) ;
    xor2 ix1124 (.Y (nx1123), .A0 (nx1125), .A1 (nx624)) ;
    xor2 ix1150 (.Y (nx1149), .A0 (nx1151), .A1 (nx1537)) ;
    xor2 ix1158 (.Y (nx1157), .A0 (nx1159), .A1 (nx274)) ;
    xor2 ix1178 (.Y (nx1177), .A0 (nx1179), .A1 (nx98)) ;
    xor2 ix1186 (.Y (nx1185), .A0 (nx1187), .A1 (nx1535)) ;
    xor2 ix945 (.Y (nx944), .A0 (nx920), .A1 (nx916)) ;
    xor2 ix943 (.Y (nx942), .A0 (nx862), .A1 (nx1541)) ;
    xor2 ix725 (.Y (nx724), .A0 (nx688), .A1 (nx1539)) ;
    xor2 ix723 (.Y (nx722), .A0 (nx628), .A1 (nx624)) ;
    xor2 ix375 (.Y (nx374), .A0 (nx338), .A1 (nx1537)) ;
    xor2 ix373 (.Y (nx372), .A0 (nx278), .A1 (nx274)) ;
    xor2 ix141 (.Y (nx140), .A0 (nx102), .A1 (nx98)) ;
    xor2 ix139 (.Y (nx138), .A0 (nx42), .A1 (nx1535)) ;
    xor2 ix1296 (.Y (nx1295), .A0 (nx1297), .A1 (nx916)) ;
    xor2 ix1307 (.Y (nx1306), .A0 (nx1308), .A1 (nx1541)) ;
    xor2 ix1318 (.Y (nx1317), .A0 (nx1319), .A1 (nx1539)) ;
    xor2 ix1323 (.Y (nx1322), .A0 (nx1324), .A1 (nx624)) ;
    xor2 ix1345 (.Y (nx1344), .A0 (nx1346), .A1 (nx1537)) ;
    xor2 ix1350 (.Y (nx1349), .A0 (nx1351), .A1 (nx274)) ;
    xor2 ix1366 (.Y (nx1365), .A0 (nx1367), .A1 (nx98)) ;
    xor2 ix1376 (.Y (nx1375), .A0 (nx1377), .A1 (nx1535)) ;
    xor2 ix1137 (.Y (nx1136), .A0 (nx928), .A1 (nx916)) ;
    xor2 ix1139 (.Y (nx1138), .A0 (nx870), .A1 (nx822)) ;
    xor2 ix705 (.Y (nx704), .A0 (nx696), .A1 (nx650)) ;
    xor2 ix703 (.Y (nx702), .A0 (nx636), .A1 (nx624)) ;
    xor2 ix355 (.Y (nx354), .A0 (nx346), .A1 (nx300)) ;
    xor2 ix353 (.Y (nx352), .A0 (nx286), .A1 (nx274)) ;
    xor2 ix121 (.Y (nx120), .A0 (nx110), .A1 (nx98)) ;
    xor2 ix119 (.Y (nx118), .A0 (nx50), .A1 (nx6)) ;
    xor2 ix1436 (.Y (nx1435), .A0 (nx6), .A1 (nx1437)) ;
    xor2 ix1449 (.Y (nx1448), .A0 (nx1450), .A1 (nx300)) ;
    xor2 ix1466 (.Y (nx1465), .A0 (nx1467), .A1 (nx650)) ;
    xor2 ix825 (.Y (nx824), .A0 (nx814), .A1 (nx822)) ;
    inv01 ix1534 (.Y (nx1535), .A (nx1189)) ;
    inv01 ix1536 (.Y (nx1537), .A (nx1153)) ;
    inv01 ix1538 (.Y (nx1539), .A (nx1119)) ;
    inv01 ix1540 (.Y (nx1541), .A (nx1099)) ;
endmodule

