-- mult_DFarch.vhd
-- Jean P. Walker
-- Architecture file using dataflow for multiplier entity.

architecture dataflow of multiplier is
begin
  C <= A * B;
end architecture;
